**** Created by MC2: Version 2010.02.00.a on 2022/02/24, 21:11:02 

************************************************************************
* AUCDL NETLIST:
* 
* LIBRARY NAME:  N65LP_SP_LEAFCELL
* TOP CELL NAME: LEAFCELLS
* VIEW NAME:     SCHEMATIC
* NETLISTED ON:  DEC 22 10:05:16 2009
************************************************************************

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MCB
* VIEW NAME:    SCHEMATIC
************************************************************************
*.BIPOLAR
*.CAPA
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA

.SUBCKT S1AHSF400W40_MIO_HD D G S B
MPCH D G S B PCH L=70N W=1.2u M=6
.ENDS

.SUBCKT S1AHSF400W40_MCB BL BLB VDDI VSSI WL
*.PININFO BL:B BLB:B VDDI:B VSSI:B WL:B
MPCHPU0 VDDI BLB_IN BL_IN VDDI PCHPU_WISR L=0.065U W=0.080U M=1
MPCHPU1 BLB_IN BL_IN VDDI VDDI PCHPU_WISR L=0.065U W=0.080U M=1
MNCHPD1 BLB_IN BL_IN VSSI VSSI NCHPD_WISR L=0.065U W=0.140U M=1
MNCHPD0 VSSI BLB_IN BL_IN VSSI NCHPD_WISR L=0.065U W=0.140U M=1
MNCHPG0 BL_IN WL BL VSSI NCHPG_WISR L=0.075U W=0.090U M=1
MNCHPG1 BLB WL BLB_IN VSSI NCHPG_WISR L=0.075U W=0.090U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    MCB_2X16_SB_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_2X16_SB_CHAR BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] 
+ BL[9] BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BLB[0] BLB[1] BLB[2] BLB[3] 
+ BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] 
+ BLB[14] BLB[15] VDDI VSSI WL[0] WL[1]
*.PININFO WL[0]:I WL[1]:I BL[0]:B BL[1]:B BL[2]:B BL[3]:B BL[4]:B BL[5]:B 
*.PININFO BL[6]:B BL[7]:B BL[8]:B BL[9]:B BL[10]:B BL[11]:B BL[12]:B BL[13]:B 
*.PININFO BL[14]:B BL[15]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B BLB[4]:B 
*.PININFO BLB[5]:B BLB[6]:B BLB[7]:B BLB[8]:B BLB[9]:B BLB[10]:B BLB[11]:B 
*.PININFO BLB[12]:B BLB[13]:B BLB[14]:B BLB[15]:B VDDI:B VSSI:B
XMCB_0<0> BL[0] BLB[0] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<1> BL[1] BLB[1] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<2> BL[2] BLB[2] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<3> BL[3] BLB[3] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<4> BL[4] BLB[4] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<5> BL[5] BLB[5] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<6> BL[6] BLB[6] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<7> BL[7] BLB[7] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<8> BL[8] BLB[8] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<9> BL[9] BLB[9] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<10> BL[10] BLB[10] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<11> BL[11] BLB[11] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<12> BL[12] BLB[12] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<13> BL[13] BLB[13] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<14> BL[14] BLB[14] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<15> BL[15] BLB[15] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_1<0> BL[0] BLB[0] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<1> BL[1] BLB[1] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<2> BL[2] BLB[2] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<3> BL[3] BLB[3] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<4> BL[4] BLB[4] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<5> BL[5] BLB[5] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<6> BL[6] BLB[6] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<7> BL[7] BLB[7] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<8> BL[8] BLB[8] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<9> BL[9] BLB[9] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<10> BL[10] BLB[10] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<11> BL[11] BLB[11] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<12> BL[12] BLB[12] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<13> BL[13] BLB[13] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<14> BL[14] BLB[14] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<15> BL[15] BLB[15] VDDI VSSI WL[1] S1AHSF400W40_MCB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    MCB_2X8_SB_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_2X8_SB_CHAR BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BLB[0] 
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] VDDI VSSI WL[0] WL[1]
*.PININFO WL[0]:I WL[1]:I BL[0]:B BL[1]:B BL[2]:B BL[3]:B BL[4]:B BL[5]:B 
*.PININFO BL[6]:B BL[7]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B BLB[4]:B 
*.PININFO BLB[5]:B BLB[6]:B BLB[7]:B VDDI:B VSSI:B
XMCB_0<0> BL[0] BLB[0] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<1> BL[1] BLB[1] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<2> BL[2] BLB[2] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<3> BL[3] BLB[3] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<4> BL[4] BLB[4] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<5> BL[5] BLB[5] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<6> BL[6] BLB[6] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<7> BL[7] BLB[7] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_1<0> BL[0] BLB[0] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<1> BL[1] BLB[1] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<2> BL[2] BLB[2] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<3> BL[3] BLB[3] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<4> BL[4] BLB[4] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<5> BL[5] BLB[5] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<6> BL[6] BLB[6] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<7> BL[7] BLB[7] VDDI VSSI WL[1] S1AHSF400W40_MCB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    MCB_2X4_SB_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_2X4_SB_CHAR BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] 
+ VDDI VSSI WL[0] WL[1]
*.PININFO WL[0]:I WL[1]:I BL[0]:B BL[1]:B BL[2]:B BL[3]:B BLB[0]:B BLB[1]:B 
*.PININFO BLB[2]:B BLB[3]:B VDDI:B VSSI:B
XMCB_0<0> BL[0] BLB[0] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<1> BL[1] BLB[1] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<2> BL[2] BLB[2] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<3> BL[3] BLB[3] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_1<0> BL[0] BLB[0] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<1> BL[1] BLB[1] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<2> BL[2] BLB[2] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<3> BL[3] BLB[3] VDDI VSSI WL[1] S1AHSF400W40_MCB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_ARR_WLLD_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_ARR_WLLD_SIM CVDDI VDDHD VDDI VSSI WL_LT[0] WL_LT[1] WL_RT[0] 
+ WL_RT[1]
*.PININFO CVDDI:B VDDHD:B VDDI:B VSSI:B WL_LT[0]:B WL_LT[1]:B WL_RT[0]:B 
*.PININFO WL_RT[1]:B
XI265 NET11[0] NET11[1] NET11[2] NET11[3] NET7[0] NET7[1] NET7[2] NET7[3] 
+ NET10 NET9 NET8[0] NET8[1] S1AHSF400W40_MCB_2X4_SB_CHAR
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    TKBL_EDGE
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TKBL_EDGE BLB_EDGE BL_EDGE CVDDI VSSI WL WL_TK TIEH
*.PININFO WL:I WL_TK:I BLB_EDGE:B BL_EDGE:B CVDDI:B VSSI:B TIEH:B
MNCHPD0 VSSI TIEH BL_TK_IN VSSI NCHPD_WISR L=0.065U W=0.140U M=1
MNCHPD1 BLB_IN BL_TK_IN VSSI VSSI NCHPD_WISR L=0.065U W=0.140U M=1
MPCHPU0 CVDDI TIEH BL_TK_IN CVDDI PCHPU_WISR L=0.065U W=0.080U M=1
MPCHPU1 TIEH BL_TK_IN CVDDI CVDDI PCHPU_WISR L=0.065U W=0.080U M=1
MNCHPG1 BLB_IN WL BLB_EDGE VSSI NCHPG_WISR L=0.075U W=0.090U M=1
MNCHPG0 BL_EDGE WL_TK BL_TK_IN VSSI NCHPG_WISR L=0.075U W=0.090U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    TKBL_BCELL
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TKBL_BCELL BLB BL_TK CVDDI VSSI WL WL_TK TIEH
*.PININFO WL:I WL_TK:I BLB:B BL_TK:B CVDDI:B VSSI:B TIEH:B
MNCHPD1 BLB_IN BL_TK_IN VSSI VSSI NCHPD_WISR L=0.065U W=0.140U M=1
MNCHPD0 VSSI TIEH BL_TK_IN VSSI NCHPD_WISR L=0.065U W=0.140U M=1
MPCHPU0 CVDDI TIEH BL_TK_IN CVDDI PCHPU_WISR L=0.065U W=0.080U M=1
MPCHPU1 TIEH BL_TK_IN CVDDI CVDDI PCHPU_WISR L=0.065U W=0.080U M=1
MNCHPG1 BLB_IN WL BLB VSSI NCHPG_WISR L=0.075U W=0.090U M=1
MNCHPG0 BL_TK WL_TK BL_TK_IN VSSI NCHPG_WISR L=0.075U W=0.090U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    TRKNOR_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TRKNOR_CHAR BLB BLB_EDGE BL_EDGE BL_TK VDDI VSSI WL WL_TK TIEH
*.PININFO WL:I WL_TK:I TIEH:I BLB:B BLB_EDGE:B BL_EDGE:B BL_TK:B VDDI:B VSSI:B
XTKBL_EDGE BLB_EDGE BL_EDGE VDDI VSSI WL WL_TK TIEH S1AHSF400W40_TKBL_EDGE
XTKBL_BCELL BLB BL_TK VDDI VSSI WL WL_TK TIEH S1AHSF400W40_TKBL_BCELL
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    TRKNORX2_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TRKNORX2_CHAR BL_TK VDDI VSSI WL[0] WL[1] WL_TK[0] WL_TK[1] FLOAT1 
+ FLOAT2 FLOAT3 FLOAT4 TIEH
*.PININFO WL[0]:I WL[1]:I WL_TK[0]:I WL_TK[1]:I TIEH:I BL_TK:B VDDI:B VSSI:B 
*.PININFO FLOAT1:B FLOAT2:B FLOAT3:B FLOAT4:B
XTRKNOR_0 FLOAT4 FLOAT1 FLOAT3 BL_TK VDDI VSSI WL[0] WL_TK[0] TIEH 
+ S1AHSF400W40_TRKNOR_CHAR
XTRKNOR_1 FLOAT4 FLOAT1 FLOAT2 BL_TK VDDI VSSI WL[1] WL_TK[1] TIEH 
+ S1AHSF400W40_TRKNOR_CHAR
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    TRKNORX4_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TRKNORX4_CHAR BL_TK VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL_TK[0] 
+ WL_TK[1] WL_TK[2] WL_TK[3] FLOAT1[0] FLOAT1[1] FLOAT2 FLOAT3 FLOAT4[0] 
+ FLOAT4[1] TIEH
*.PININFO WL[0]:I WL[1]:I WL[2]:I WL[3]:I WL_TK[0]:I WL_TK[1]:I WL_TK[2]:I 
*.PININFO WL_TK[3]:I TIEH:I BL_TK:B VDDI:B VSSI:B FLOAT1[0]:B FLOAT1[1]:B 
*.PININFO FLOAT2:B FLOAT3:B FLOAT4[0]:B FLOAT4[1]:B
XTRKNORX2_0 BL_TK VDDI VSSI WL[0] WL[1] WL_TK[0] WL_TK[1] FLOAT1[0] NET30 
+ FLOAT3 FLOAT4[0] TIEH S1AHSF400W40_TRKNORX2_CHAR
XTRKNORX2_1 BL_TK VDDI VSSI WL[2] WL[3] WL_TK[2] WL_TK[3] FLOAT1[1] FLOAT2 
+ NET30 FLOAT4[1] TIEH S1AHSF400W40_TRKNORX2_CHAR
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    TRKNORX16_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TRKNORX16_CHAR BL_TK VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL_TK[0] 
+ WL_TK[1] WL_TK[2] WL_TK[3] WL_TK[4] WL_TK[5] WL_TK[6] WL_TK[7] WL_TK[8] 
+ WL_TK[9] WL_TK[10] WL_TK[11] WL_TK[12] WL_TK[13] WL_TK[14] WL_TK[15] 
+ FLOAT1[0] FLOAT1[1] FLOAT1[2] FLOAT1[3] FLOAT1[4] FLOAT1[5] FLOAT1[6] 
+ FLOAT1[7] FLOAT2 FLOAT3 FLOAT4[0] FLOAT4[1] FLOAT4[2] FLOAT4[3] FLOAT4[4] 
+ FLOAT4[5] FLOAT4[6] FLOAT4[7] TIEH
*.PININFO WL[0]:I WL[1]:I WL[2]:I WL[3]:I WL[4]:I WL[5]:I WL[6]:I WL[7]:I 
*.PININFO WL[8]:I WL[9]:I WL[10]:I WL[11]:I WL[12]:I WL[13]:I WL[14]:I 
*.PININFO WL[15]:I WL_TK[0]:I WL_TK[1]:I WL_TK[2]:I WL_TK[3]:I WL_TK[4]:I 
*.PININFO WL_TK[5]:I WL_TK[6]:I WL_TK[7]:I WL_TK[8]:I WL_TK[9]:I WL_TK[10]:I 
*.PININFO WL_TK[11]:I WL_TK[12]:I WL_TK[13]:I WL_TK[14]:I WL_TK[15]:I BL_TK:B 
*.PININFO VDDI:B VSSI:B FLOAT1[0]:B FLOAT1[1]:B FLOAT1[2]:B FLOAT1[3]:B 
*.PININFO FLOAT1[4]:B FLOAT1[5]:B FLOAT1[6]:B FLOAT1[7]:B FLOAT2:B FLOAT3:B 
*.PININFO FLOAT4[0]:B FLOAT4[1]:B FLOAT4[2]:B FLOAT4[3]:B FLOAT4[4]:B 
*.PININFO FLOAT4[5]:B FLOAT4[6]:B FLOAT4[7]:B TIEH:B
XTRKNORX4_2 BL_TK VDDI VSSI WL[8] WL[9] WL[10] WL[11] WL_TK[8] WL_TK[9] 
+ WL_TK[10] WL_TK[11] FLOAT1[4] FLOAT1[5] NET29 NET39 FLOAT4[4] FLOAT4[5] TIEH 
+ S1AHSF400W40_TRKNORX4_CHAR
XTRKNORX4_1 BL_TK VDDI VSSI WL[4] WL[5] WL[6] WL[7] WL_TK[4] WL_TK[5] WL_TK[6] 
+ WL_TK[7] FLOAT1[2] FLOAT1[3] NET39 NET49 FLOAT4[2] FLOAT4[3] TIEH 
+ S1AHSF400W40_TRKNORX4_CHAR
XTRKNORX4_3 BL_TK VDDI VSSI WL[12] WL[13] WL[14] WL[15] WL_TK[12] WL_TK[13] 
+ WL_TK[14] WL_TK[15] FLOAT1[6] FLOAT1[7] FLOAT2 NET29 FLOAT4[6] FLOAT4[7] 
+ TIEH S1AHSF400W40_TRKNORX4_CHAR
XTRKNORX4_0 BL_TK VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL_TK[0] WL_TK[1] WL_TK[2] 
+ WL_TK[3] FLOAT1[0] FLOAT1[1] NET49 FLOAT3 FLOAT4[0] FLOAT4[1] TIEH 
+ S1AHSF400W40_TRKNORX4_CHAR
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    TRKNORX64_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TRKNORX64_CHAR BL_TK VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL_TK[0] WL_TK[1] WL_TK[2] WL_TK[3] WL_TK[4] WL_TK[5] 
+ WL_TK[6] WL_TK[7] WL_TK[8] WL_TK[9] WL_TK[10] WL_TK[11] WL_TK[12] WL_TK[13] 
+ WL_TK[14] WL_TK[15] WL_TK[16] WL_TK[17] WL_TK[18] WL_TK[19] WL_TK[20] 
+ WL_TK[21] WL_TK[22] WL_TK[23] WL_TK[24] WL_TK[25] WL_TK[26] WL_TK[27] 
+ WL_TK[28] WL_TK[29] WL_TK[30] WL_TK[31] WL_TK[32] WL_TK[33] WL_TK[34] 
+ WL_TK[35] WL_TK[36] WL_TK[37] WL_TK[38] WL_TK[39] WL_TK[40] WL_TK[41] 
+ WL_TK[42] WL_TK[43] WL_TK[44] WL_TK[45] WL_TK[46] WL_TK[47] WL_TK[48] 
+ WL_TK[49] WL_TK[50] WL_TK[51] WL_TK[52] WL_TK[53] WL_TK[54] WL_TK[55] 
+ WL_TK[56] WL_TK[57] WL_TK[58] WL_TK[59] WL_TK[60] WL_TK[61] WL_TK[62] 
+ WL_TK[63] FLOAT1[31] FLOAT1[30] FLOAT1[29] FLOAT1[28] FLOAT1[27] FLOAT1[26] 
+ FLOAT1[25] FLOAT1[24] FLOAT1[23] FLOAT1[22] FLOAT1[21] FLOAT1[20] FLOAT1[19] 
+ FLOAT1[18] FLOAT1[17] FLOAT1[16] FLOAT1[15] FLOAT1[14] FLOAT1[13] FLOAT1[12] 
+ FLOAT1[11] FLOAT1[10] FLOAT1[9] FLOAT1[8] FLOAT1[7] FLOAT1[6] FLOAT1[5] 
+ FLOAT1[4] FLOAT1[3] FLOAT1[2] FLOAT1[1] FLOAT1[0] FLOAT2 FLOAT3 FLOAT4[31] 
+ FLOAT4[30] FLOAT4[29] FLOAT4[28] FLOAT4[27] FLOAT4[26] FLOAT4[25] FLOAT4[24] 
+ FLOAT4[23] FLOAT4[22] FLOAT4[21] FLOAT4[20] FLOAT4[19] FLOAT4[18] FLOAT4[17] 
+ FLOAT4[16] FLOAT4[15] FLOAT4[14] FLOAT4[13] FLOAT4[12] FLOAT4[11] FLOAT4[10] 
+ FLOAT4[9] FLOAT4[8] FLOAT4[7] FLOAT4[6] FLOAT4[5] FLOAT4[4] FLOAT4[3] 
+ FLOAT4[2] FLOAT4[1] FLOAT4[0] TIEH
*.PININFO WL[0]:I WL[1]:I WL[2]:I WL[3]:I WL[4]:I WL[5]:I WL[6]:I WL[7]:I 
*.PININFO WL[8]:I WL[9]:I WL[10]:I WL[11]:I WL[12]:I WL[13]:I WL[14]:I 
*.PININFO WL[15]:I WL[16]:I WL[17]:I WL[18]:I WL[19]:I WL[20]:I WL[21]:I 
*.PININFO WL[22]:I WL[23]:I WL[24]:I WL[25]:I WL[26]:I WL[27]:I WL[28]:I 
*.PININFO WL[29]:I WL[30]:I WL[31]:I WL[32]:I WL[33]:I WL[34]:I WL[35]:I 
*.PININFO WL[36]:I WL[37]:I WL[38]:I WL[39]:I WL[40]:I WL[41]:I WL[42]:I 
*.PININFO WL[43]:I WL[44]:I WL[45]:I WL[46]:I WL[47]:I WL[48]:I WL[49]:I 
*.PININFO WL[50]:I WL[51]:I WL[52]:I WL[53]:I WL[54]:I WL[55]:I WL[56]:I 
*.PININFO WL[57]:I WL[58]:I WL[59]:I WL[60]:I WL[61]:I WL[62]:I WL[63]:I 
*.PININFO WL_TK[0]:I WL_TK[1]:I WL_TK[2]:I WL_TK[3]:I WL_TK[4]:I WL_TK[5]:I 
*.PININFO WL_TK[6]:I WL_TK[7]:I WL_TK[8]:I WL_TK[9]:I WL_TK[10]:I WL_TK[11]:I 
*.PININFO WL_TK[12]:I WL_TK[13]:I WL_TK[14]:I WL_TK[15]:I WL_TK[16]:I 
*.PININFO WL_TK[17]:I WL_TK[18]:I WL_TK[19]:I WL_TK[20]:I WL_TK[21]:I 
*.PININFO WL_TK[22]:I WL_TK[23]:I WL_TK[24]:I WL_TK[25]:I WL_TK[26]:I 
*.PININFO WL_TK[27]:I WL_TK[28]:I WL_TK[29]:I WL_TK[30]:I WL_TK[31]:I 
*.PININFO WL_TK[32]:I WL_TK[33]:I WL_TK[34]:I WL_TK[35]:I WL_TK[36]:I 
*.PININFO WL_TK[37]:I WL_TK[38]:I WL_TK[39]:I WL_TK[40]:I WL_TK[41]:I 
*.PININFO WL_TK[42]:I WL_TK[43]:I WL_TK[44]:I WL_TK[45]:I WL_TK[46]:I 
*.PININFO WL_TK[47]:I WL_TK[48]:I WL_TK[49]:I WL_TK[50]:I WL_TK[51]:I 
*.PININFO WL_TK[52]:I WL_TK[53]:I WL_TK[54]:I WL_TK[55]:I WL_TK[56]:I 
*.PININFO WL_TK[57]:I WL_TK[58]:I WL_TK[59]:I WL_TK[60]:I WL_TK[61]:I 
*.PININFO WL_TK[62]:I WL_TK[63]:I BL_TK:B VDDI:B VSSI:B FLOAT1[31]:B 
*.PININFO FLOAT1[30]:B FLOAT1[29]:B FLOAT1[28]:B FLOAT1[27]:B FLOAT1[26]:B 
*.PININFO FLOAT1[25]:B FLOAT1[24]:B FLOAT1[23]:B FLOAT1[22]:B FLOAT1[21]:B 
*.PININFO FLOAT1[20]:B FLOAT1[19]:B FLOAT1[18]:B FLOAT1[17]:B FLOAT1[16]:B 
*.PININFO FLOAT1[15]:B FLOAT1[14]:B FLOAT1[13]:B FLOAT1[12]:B FLOAT1[11]:B 
*.PININFO FLOAT1[10]:B FLOAT1[9]:B FLOAT1[8]:B FLOAT1[7]:B FLOAT1[6]:B 
*.PININFO FLOAT1[5]:B FLOAT1[4]:B FLOAT1[3]:B FLOAT1[2]:B FLOAT1[1]:B 
*.PININFO FLOAT1[0]:B FLOAT2:B FLOAT3:B FLOAT4[31]:B FLOAT4[30]:B FLOAT4[29]:B 
*.PININFO FLOAT4[28]:B FLOAT4[27]:B FLOAT4[26]:B FLOAT4[25]:B FLOAT4[24]:B 
*.PININFO FLOAT4[23]:B FLOAT4[22]:B FLOAT4[21]:B FLOAT4[20]:B FLOAT4[19]:B 
*.PININFO FLOAT4[18]:B FLOAT4[17]:B FLOAT4[16]:B FLOAT4[15]:B FLOAT4[14]:B 
*.PININFO FLOAT4[13]:B FLOAT4[12]:B FLOAT4[11]:B FLOAT4[10]:B FLOAT4[9]:B 
*.PININFO FLOAT4[8]:B FLOAT4[7]:B FLOAT4[6]:B FLOAT4[5]:B FLOAT4[4]:B 
*.PININFO FLOAT4[3]:B FLOAT4[2]:B FLOAT4[1]:B FLOAT4[0]:B TIEH:B
XTRKNORX16_3 BL_TK VDDI VSSI WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] 
+ WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] WL_TK[48] 
+ WL_TK[49] WL_TK[50] WL_TK[51] WL_TK[52] WL_TK[53] WL_TK[54] WL_TK[55] 
+ WL_TK[56] WL_TK[57] WL_TK[58] WL_TK[59] WL_TK[60] WL_TK[61] WL_TK[62] 
+ WL_TK[63] FLOAT1[24] FLOAT1[25] FLOAT1[26] FLOAT1[27] FLOAT1[28] FLOAT1[29] 
+ FLOAT1[30] FLOAT1[31] FLOAT2 NET26 FLOAT4[24] FLOAT4[25] FLOAT4[26] 
+ FLOAT4[27] FLOAT4[28] FLOAT4[29] FLOAT4[30] FLOAT4[31] TIEH S1AHSF400W40_TRKNORX16_CHAR
XTRKNORX16_2 BL_TK VDDI VSSI WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL_TK[32] 
+ WL_TK[33] WL_TK[34] WL_TK[35] WL_TK[36] WL_TK[37] WL_TK[38] WL_TK[39] 
+ WL_TK[40] WL_TK[41] WL_TK[42] WL_TK[43] WL_TK[44] WL_TK[45] WL_TK[46] 
+ WL_TK[47] FLOAT1[16] FLOAT1[17] FLOAT1[18] FLOAT1[19] FLOAT1[20] FLOAT1[21] 
+ FLOAT1[22] FLOAT1[23] NET26 NET36 FLOAT4[16] FLOAT4[17] FLOAT4[18] 
+ FLOAT4[19] FLOAT4[20] FLOAT4[21] FLOAT4[22] FLOAT4[23] TIEH S1AHSF400W40_TRKNORX16_CHAR
XTRKNORX16_1 BL_TK VDDI VSSI WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] 
+ WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL_TK[16] 
+ WL_TK[17] WL_TK[18] WL_TK[19] WL_TK[20] WL_TK[21] WL_TK[22] WL_TK[23] 
+ WL_TK[24] WL_TK[25] WL_TK[26] WL_TK[27] WL_TK[28] WL_TK[29] WL_TK[30] 
+ WL_TK[31] FLOAT1[8] FLOAT1[9] FLOAT1[10] FLOAT1[11] FLOAT1[12] FLOAT1[13] 
+ FLOAT1[14] FLOAT1[15] NET36 NET47 FLOAT4[8] FLOAT4[9] FLOAT4[10] FLOAT4[11] 
+ FLOAT4[12] FLOAT4[13] FLOAT4[14] FLOAT4[15] TIEH S1AHSF400W40_TRKNORX16_CHAR
XTRKNORX16_0 BL_TK VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] 
+ WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL_TK[0] WL_TK[1] 
+ WL_TK[2] WL_TK[3] WL_TK[4] WL_TK[5] WL_TK[6] WL_TK[7] WL_TK[8] WL_TK[9] 
+ WL_TK[10] WL_TK[11] WL_TK[12] WL_TK[13] WL_TK[14] WL_TK[15] FLOAT1[0] 
+ FLOAT1[1] FLOAT1[2] FLOAT1[3] FLOAT1[4] FLOAT1[5] FLOAT1[6] FLOAT1[7] NET47 
+ FLOAT3 FLOAT4[0] FLOAT4[1] FLOAT4[2] FLOAT4[3] FLOAT4[4] FLOAT4[5] FLOAT4[6] 
+ FLOAT4[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    TKBL_S384_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TKBL_S384_CHAR BL_TK VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] WL_TK[0] WL_TK[1] WL_TK[2] WL_TK[3] WL_TK[4] 
+ WL_TK[5] WL_TK[6] WL_TK[7] WL_TK[8] WL_TK[9] WL_TK[10] WL_TK[11] WL_TK[12] 
+ WL_TK[13] WL_TK[14] WL_TK[15] WL_TK[16] WL_TK[17] WL_TK[18] WL_TK[19] 
+ WL_TK[20] WL_TK[21] WL_TK[22] WL_TK[23] WL_TK[24] WL_TK[25] WL_TK[26] 
+ WL_TK[27] WL_TK[28] WL_TK[29] WL_TK[30] WL_TK[31] WL_TK[32] WL_TK[33] 
+ WL_TK[34] WL_TK[35] WL_TK[36] WL_TK[37] WL_TK[38] WL_TK[39] WL_TK[40] 
+ WL_TK[41] WL_TK[42] WL_TK[43] WL_TK[44] WL_TK[45] WL_TK[46] WL_TK[47] 
+ WL_TK[48] WL_TK[49] WL_TK[50] WL_TK[51] WL_TK[52] WL_TK[53] WL_TK[54] 
+ WL_TK[55] WL_TK[56] WL_TK[57] WL_TK[58] WL_TK[59] WL_TK[60] WL_TK[61] 
+ WL_TK[62] WL_TK[63] WL_TK[64] WL_TK[65] WL_TK[66] WL_TK[67] WL_TK[68] 
+ WL_TK[69] WL_TK[70] WL_TK[71] WL_TK[72] WL_TK[73] WL_TK[74] WL_TK[75] 
+ WL_TK[76] WL_TK[77] WL_TK[78] WL_TK[79] WL_TK[80] WL_TK[81] WL_TK[82] 
+ WL_TK[83] WL_TK[84] WL_TK[85] WL_TK[86] WL_TK[87] WL_TK[88] WL_TK[89] 
+ WL_TK[90] WL_TK[91] WL_TK[92] WL_TK[93] WL_TK[94] WL_TK[95] WL_TK[96] 
+ WL_TK[97] WL_TK[98] WL_TK[99] WL_TK[100] WL_TK[101] WL_TK[102] WL_TK[103] 
+ WL_TK[104] WL_TK[105] WL_TK[106] WL_TK[107] WL_TK[108] WL_TK[109] WL_TK[110] 
+ WL_TK[111] WL_TK[112] WL_TK[113] WL_TK[114] WL_TK[115] WL_TK[116] WL_TK[117] 
+ WL_TK[118] WL_TK[119] WL_TK[120] WL_TK[121] WL_TK[122] WL_TK[123] WL_TK[124] 
+ WL_TK[125] WL_TK[126] WL_TK[127] WL_TK[128] WL_TK[129] WL_TK[130] WL_TK[131] 
+ WL_TK[132] WL_TK[133] WL_TK[134] WL_TK[135] WL_TK[136] WL_TK[137] WL_TK[138] 
+ WL_TK[139] WL_TK[140] WL_TK[141] WL_TK[142] WL_TK[143] WL_TK[144] WL_TK[145] 
+ WL_TK[146] WL_TK[147] WL_TK[148] WL_TK[149] WL_TK[150] WL_TK[151] WL_TK[152] 
+ WL_TK[153] WL_TK[154] WL_TK[155] WL_TK[156] WL_TK[157] WL_TK[158] WL_TK[159] 
+ WL_TK[160] WL_TK[161] WL_TK[162] WL_TK[163] WL_TK[164] WL_TK[165] WL_TK[166] 
+ WL_TK[167] WL_TK[168] WL_TK[169] WL_TK[170] WL_TK[171] WL_TK[172] WL_TK[173] 
+ WL_TK[174] WL_TK[175] WL_TK[176] WL_TK[177] WL_TK[178] WL_TK[179] WL_TK[180] 
+ WL_TK[181] WL_TK[182] WL_TK[183] WL_TK[184] WL_TK[185] WL_TK[186] WL_TK[187] 
+ WL_TK[188] WL_TK[189] WL_TK[190] WL_TK[191] WL_TK[192] WL_TK[193] WL_TK[194] 
+ WL_TK[195] WL_TK[196] WL_TK[197] WL_TK[198] WL_TK[199] WL_TK[200] WL_TK[201] 
+ WL_TK[202] WL_TK[203] WL_TK[204] WL_TK[205] WL_TK[206] WL_TK[207] WL_TK[208] 
+ WL_TK[209] WL_TK[210] WL_TK[211] WL_TK[212] WL_TK[213] WL_TK[214] WL_TK[215] 
+ WL_TK[216] WL_TK[217] WL_TK[218] WL_TK[219] WL_TK[220] WL_TK[221] WL_TK[222] 
+ WL_TK[223] WL_TK[224] WL_TK[225] WL_TK[226] WL_TK[227] WL_TK[228] WL_TK[229] 
+ WL_TK[230] WL_TK[231] WL_TK[232] WL_TK[233] WL_TK[234] WL_TK[235] WL_TK[236] 
+ WL_TK[237] WL_TK[238] WL_TK[239] WL_TK[240] WL_TK[241] WL_TK[242] WL_TK[243] 
+ WL_TK[244] WL_TK[245] WL_TK[246] WL_TK[247] WL_TK[248] WL_TK[249] WL_TK[250] 
+ WL_TK[251] WL_TK[252] WL_TK[253] WL_TK[254] WL_TK[255] WL_TK[256] WL_TK[257] 
+ WL_TK[258] WL_TK[259] WL_TK[260] WL_TK[261] WL_TK[262] WL_TK[263] WL_TK[264] 
+ WL_TK[265] WL_TK[266] WL_TK[267] WL_TK[268] WL_TK[269] WL_TK[270] WL_TK[271] 
+ WL_TK[272] WL_TK[273] WL_TK[274] WL_TK[275] WL_TK[276] WL_TK[277] WL_TK[278] 
+ WL_TK[279] WL_TK[280] WL_TK[281] WL_TK[282] WL_TK[283] WL_TK[284] WL_TK[285] 
+ WL_TK[286] WL_TK[287] WL_TK[288] WL_TK[289] WL_TK[290] WL_TK[291] WL_TK[292] 
+ WL_TK[293] WL_TK[294] WL_TK[295] WL_TK[296] WL_TK[297] WL_TK[298] WL_TK[299] 
+ WL_TK[300] WL_TK[301] WL_TK[302] WL_TK[303] WL_TK[304] WL_TK[305] WL_TK[306] 
+ WL_TK[307] WL_TK[308] WL_TK[309] WL_TK[310] WL_TK[311] WL_TK[312] WL_TK[313] 
+ WL_TK[314] WL_TK[315] WL_TK[316] WL_TK[317] WL_TK[318] WL_TK[319] WL_TK[320] 
+ WL_TK[321] WL_TK[322] WL_TK[323] WL_TK[324] WL_TK[325] WL_TK[326] WL_TK[327] 
+ WL_TK[328] WL_TK[329] WL_TK[330] WL_TK[331] WL_TK[332] WL_TK[333] WL_TK[334] 
+ WL_TK[335] WL_TK[336] WL_TK[337] WL_TK[338] WL_TK[339] WL_TK[340] WL_TK[341] 
+ WL_TK[342] WL_TK[343] WL_TK[344] WL_TK[345] WL_TK[346] WL_TK[347] WL_TK[348] 
+ WL_TK[349] WL_TK[350] WL_TK[351] WL_TK[352] WL_TK[353] WL_TK[354] WL_TK[355] 
+ WL_TK[356] WL_TK[357] WL_TK[358] WL_TK[359] WL_TK[360] WL_TK[361] WL_TK[362] 
+ WL_TK[363] WL_TK[364] WL_TK[365] WL_TK[366] WL_TK[367] WL_TK[368] WL_TK[369] 
+ WL_TK[370] WL_TK[371] WL_TK[372] WL_TK[373] WL_TK[374] WL_TK[375] WL_TK[376] 
+ WL_TK[377] WL_TK[378] WL_TK[379] WL_TK[380] WL_TK[381] WL_TK[382] WL_TK[383] 
+ WL_TK[384] WL_TK[385] WL_TK[386] WL_TK[387] WL_TK[388] WL_TK[389] WL_TK[390] 
+ WL_TK[391] WL_TK[392] WL_TK[393] WL_TK[394] WL_TK[395] WL_TK[396] WL_TK[397] 
+ WL_TK[398] WL_TK[399] WL_TK[400] WL_TK[401] WL_TK[402] WL_TK[403] WL_TK[404] 
+ WL_TK[405] WL_TK[406] WL_TK[407] WL_TK[408] WL_TK[409] WL_TK[410] WL_TK[411] 
+ WL_TK[412] WL_TK[413] WL_TK[414] WL_TK[415] WL_TK[416] WL_TK[417] WL_TK[418] 
+ WL_TK[419] WL_TK[420] WL_TK[421] WL_TK[422] WL_TK[423] WL_TK[424] WL_TK[425] 
+ WL_TK[426] WL_TK[427] WL_TK[428] WL_TK[429] WL_TK[430] WL_TK[431] WL_TK[432] 
+ WL_TK[433] WL_TK[434] WL_TK[435] WL_TK[436] WL_TK[437] WL_TK[438] WL_TK[439] 
+ WL_TK[440] WL_TK[441] WL_TK[442] WL_TK[443] WL_TK[444] WL_TK[445] WL_TK[446] 
+ WL_TK[447] WL_TK[448] WL_TK[449] WL_TK[450] WL_TK[451] WL_TK[452] WL_TK[453] 
+ WL_TK[454] WL_TK[455] WL_TK[456] WL_TK[457] WL_TK[458] WL_TK[459] WL_TK[460] 
+ WL_TK[461] WL_TK[462] WL_TK[463] WL_TK[464] WL_TK[465] WL_TK[466] WL_TK[467] 
+ WL_TK[468] WL_TK[469] WL_TK[470] WL_TK[471] WL_TK[472] WL_TK[473] WL_TK[474] 
+ WL_TK[475] WL_TK[476] WL_TK[477] WL_TK[478] WL_TK[479] WL_TK[480] WL_TK[481] 
+ WL_TK[482] WL_TK[483] WL_TK[484] WL_TK[485] WL_TK[486] WL_TK[487] WL_TK[488] 
+ WL_TK[489] WL_TK[490] WL_TK[491] WL_TK[492] WL_TK[493] WL_TK[494] WL_TK[495] 
+ WL_TK[496] WL_TK[497] WL_TK[498] WL_TK[499] WL_TK[500] WL_TK[501] WL_TK[502] 
+ WL_TK[503] WL_TK[504] WL_TK[505] WL_TK[506] WL_TK[507] WL_TK[508] WL_TK[509] 
+ WL_TK[510] WL_TK[511] TIEH TIEL
*.PININFO BL_TK:B VDDI:B VSSI:B WL[0]:B WL[1]:B WL[2]:B WL[3]:B WL[4]:B 
*.PININFO WL[5]:B WL[6]:B WL[7]:B WL[8]:B WL[9]:B WL[10]:B WL[11]:B WL[12]:B 
*.PININFO WL[13]:B WL[14]:B WL[15]:B WL[16]:B WL[17]:B WL[18]:B WL[19]:B 
*.PININFO WL[20]:B WL[21]:B WL[22]:B WL[23]:B WL[24]:B WL[25]:B WL[26]:B 
*.PININFO WL[27]:B WL[28]:B WL[29]:B WL[30]:B WL[31]:B WL[32]:B WL[33]:B 
*.PININFO WL[34]:B WL[35]:B WL[36]:B WL[37]:B WL[38]:B WL[39]:B WL[40]:B 
*.PININFO WL[41]:B WL[42]:B WL[43]:B WL[44]:B WL[45]:B WL[46]:B WL[47]:B 
*.PININFO WL[48]:B WL[49]:B WL[50]:B WL[51]:B WL[52]:B WL[53]:B WL[54]:B 
*.PININFO WL[55]:B WL[56]:B WL[57]:B WL[58]:B WL[59]:B WL[60]:B WL[61]:B 
*.PININFO WL[62]:B WL[63]:B WL[64]:B WL[65]:B WL[66]:B WL[67]:B WL[68]:B 
*.PININFO WL[69]:B WL[70]:B WL[71]:B WL[72]:B WL[73]:B WL[74]:B WL[75]:B 
*.PININFO WL[76]:B WL[77]:B WL[78]:B WL[79]:B WL[80]:B WL[81]:B WL[82]:B 
*.PININFO WL[83]:B WL[84]:B WL[85]:B WL[86]:B WL[87]:B WL[88]:B WL[89]:B 
*.PININFO WL[90]:B WL[91]:B WL[92]:B WL[93]:B WL[94]:B WL[95]:B WL[96]:B 
*.PININFO WL[97]:B WL[98]:B WL[99]:B WL[100]:B WL[101]:B WL[102]:B WL[103]:B 
*.PININFO WL[104]:B WL[105]:B WL[106]:B WL[107]:B WL[108]:B WL[109]:B 
*.PININFO WL[110]:B WL[111]:B WL[112]:B WL[113]:B WL[114]:B WL[115]:B 
*.PININFO WL[116]:B WL[117]:B WL[118]:B WL[119]:B WL[120]:B WL[121]:B 
*.PININFO WL[122]:B WL[123]:B WL[124]:B WL[125]:B WL[126]:B WL[127]:B 
*.PININFO WL[128]:B WL[129]:B WL[130]:B WL[131]:B WL[132]:B WL[133]:B 
*.PININFO WL[134]:B WL[135]:B WL[136]:B WL[137]:B WL[138]:B WL[139]:B 
*.PININFO WL[140]:B WL[141]:B WL[142]:B WL[143]:B WL[144]:B WL[145]:B 
*.PININFO WL[146]:B WL[147]:B WL[148]:B WL[149]:B WL[150]:B WL[151]:B 
*.PININFO WL[152]:B WL[153]:B WL[154]:B WL[155]:B WL[156]:B WL[157]:B 
*.PININFO WL[158]:B WL[159]:B WL[160]:B WL[161]:B WL[162]:B WL[163]:B 
*.PININFO WL[164]:B WL[165]:B WL[166]:B WL[167]:B WL[168]:B WL[169]:B 
*.PININFO WL[170]:B WL[171]:B WL[172]:B WL[173]:B WL[174]:B WL[175]:B 
*.PININFO WL[176]:B WL[177]:B WL[178]:B WL[179]:B WL[180]:B WL[181]:B 
*.PININFO WL[182]:B WL[183]:B WL[184]:B WL[185]:B WL[186]:B WL[187]:B 
*.PININFO WL[188]:B WL[189]:B WL[190]:B WL[191]:B WL[192]:B WL[193]:B 
*.PININFO WL[194]:B WL[195]:B WL[196]:B WL[197]:B WL[198]:B WL[199]:B 
*.PININFO WL[200]:B WL[201]:B WL[202]:B WL[203]:B WL[204]:B WL[205]:B 
*.PININFO WL[206]:B WL[207]:B WL[208]:B WL[209]:B WL[210]:B WL[211]:B 
*.PININFO WL[212]:B WL[213]:B WL[214]:B WL[215]:B WL[216]:B WL[217]:B 
*.PININFO WL[218]:B WL[219]:B WL[220]:B WL[221]:B WL[222]:B WL[223]:B 
*.PININFO WL[224]:B WL[225]:B WL[226]:B WL[227]:B WL[228]:B WL[229]:B 
*.PININFO WL[230]:B WL[231]:B WL[232]:B WL[233]:B WL[234]:B WL[235]:B 
*.PININFO WL[236]:B WL[237]:B WL[238]:B WL[239]:B WL[240]:B WL[241]:B 
*.PININFO WL[242]:B WL[243]:B WL[244]:B WL[245]:B WL[246]:B WL[247]:B 
*.PININFO WL[248]:B WL[249]:B WL[250]:B WL[251]:B WL[252]:B WL[253]:B 
*.PININFO WL[254]:B WL[255]:B WL[256]:B WL[257]:B WL[258]:B WL[259]:B 
*.PININFO WL[260]:B WL[261]:B WL[262]:B WL[263]:B WL[264]:B WL[265]:B 
*.PININFO WL[266]:B WL[267]:B WL[268]:B WL[269]:B WL[270]:B WL[271]:B 
*.PININFO WL[272]:B WL[273]:B WL[274]:B WL[275]:B WL[276]:B WL[277]:B 
*.PININFO WL[278]:B WL[279]:B WL[280]:B WL[281]:B WL[282]:B WL[283]:B 
*.PININFO WL[284]:B WL[285]:B WL[286]:B WL[287]:B WL[288]:B WL[289]:B 
*.PININFO WL[290]:B WL[291]:B WL[292]:B WL[293]:B WL[294]:B WL[295]:B 
*.PININFO WL[296]:B WL[297]:B WL[298]:B WL[299]:B WL[300]:B WL[301]:B 
*.PININFO WL[302]:B WL[303]:B WL[304]:B WL[305]:B WL[306]:B WL[307]:B 
*.PININFO WL[308]:B WL[309]:B WL[310]:B WL[311]:B WL[312]:B WL[313]:B 
*.PININFO WL[314]:B WL[315]:B WL[316]:B WL[317]:B WL[318]:B WL[319]:B 
*.PININFO WL[320]:B WL[321]:B WL[322]:B WL[323]:B WL[324]:B WL[325]:B 
*.PININFO WL[326]:B WL[327]:B WL[328]:B WL[329]:B WL[330]:B WL[331]:B 
*.PININFO WL[332]:B WL[333]:B WL[334]:B WL[335]:B WL[336]:B WL[337]:B 
*.PININFO WL[338]:B WL[339]:B WL[340]:B WL[341]:B WL[342]:B WL[343]:B 
*.PININFO WL[344]:B WL[345]:B WL[346]:B WL[347]:B WL[348]:B WL[349]:B 
*.PININFO WL[350]:B WL[351]:B WL[352]:B WL[353]:B WL[354]:B WL[355]:B 
*.PININFO WL[356]:B WL[357]:B WL[358]:B WL[359]:B WL[360]:B WL[361]:B 
*.PININFO WL[362]:B WL[363]:B WL[364]:B WL[365]:B WL[366]:B WL[367]:B 
*.PININFO WL[368]:B WL[369]:B WL[370]:B WL[371]:B WL[372]:B WL[373]:B 
*.PININFO WL[374]:B WL[375]:B WL[376]:B WL[377]:B WL[378]:B WL[379]:B 
*.PININFO WL[380]:B WL[381]:B WL[382]:B WL[383]:B WL[384]:B WL[385]:B 
*.PININFO WL[386]:B WL[387]:B WL[388]:B WL[389]:B WL[390]:B WL[391]:B 
*.PININFO WL[392]:B WL[393]:B WL[394]:B WL[395]:B WL[396]:B WL[397]:B 
*.PININFO WL[398]:B WL[399]:B WL[400]:B WL[401]:B WL[402]:B WL[403]:B 
*.PININFO WL[404]:B WL[405]:B WL[406]:B WL[407]:B WL[408]:B WL[409]:B 
*.PININFO WL[410]:B WL[411]:B WL[412]:B WL[413]:B WL[414]:B WL[415]:B 
*.PININFO WL[416]:B WL[417]:B WL[418]:B WL[419]:B WL[420]:B WL[421]:B 
*.PININFO WL[422]:B WL[423]:B WL[424]:B WL[425]:B WL[426]:B WL[427]:B 
*.PININFO WL[428]:B WL[429]:B WL[430]:B WL[431]:B WL[432]:B WL[433]:B 
*.PININFO WL[434]:B WL[435]:B WL[436]:B WL[437]:B WL[438]:B WL[439]:B 
*.PININFO WL[440]:B WL[441]:B WL[442]:B WL[443]:B WL[444]:B WL[445]:B 
*.PININFO WL[446]:B WL[447]:B WL[448]:B WL[449]:B WL[450]:B WL[451]:B 
*.PININFO WL[452]:B WL[453]:B WL[454]:B WL[455]:B WL[456]:B WL[457]:B 
*.PININFO WL[458]:B WL[459]:B WL[460]:B WL[461]:B WL[462]:B WL[463]:B 
*.PININFO WL[464]:B WL[465]:B WL[466]:B WL[467]:B WL[468]:B WL[469]:B 
*.PININFO WL[470]:B WL[471]:B WL[472]:B WL[473]:B WL[474]:B WL[475]:B 
*.PININFO WL[476]:B WL[477]:B WL[478]:B WL[479]:B WL[480]:B WL[481]:B 
*.PININFO WL[482]:B WL[483]:B WL[484]:B WL[485]:B WL[486]:B WL[487]:B 
*.PININFO WL[488]:B WL[489]:B WL[490]:B WL[491]:B WL[492]:B WL[493]:B 
*.PININFO WL[494]:B WL[495]:B WL[496]:B WL[497]:B WL[498]:B WL[499]:B 
*.PININFO WL[500]:B WL[501]:B WL[502]:B WL[503]:B WL[504]:B WL[505]:B 
*.PININFO WL[506]:B WL[507]:B WL[508]:B WL[509]:B WL[510]:B WL[511]:B 
*.PININFO WL_TK[0]:B WL_TK[1]:B WL_TK[2]:B WL_TK[3]:B WL_TK[4]:B WL_TK[5]:B 
*.PININFO WL_TK[6]:B WL_TK[7]:B WL_TK[8]:B WL_TK[9]:B WL_TK[10]:B WL_TK[11]:B 
*.PININFO WL_TK[12]:B WL_TK[13]:B WL_TK[14]:B WL_TK[15]:B WL_TK[16]:B 
*.PININFO WL_TK[17]:B WL_TK[18]:B WL_TK[19]:B WL_TK[20]:B WL_TK[21]:B 
*.PININFO WL_TK[22]:B WL_TK[23]:B WL_TK[24]:B WL_TK[25]:B WL_TK[26]:B 
*.PININFO WL_TK[27]:B WL_TK[28]:B WL_TK[29]:B WL_TK[30]:B WL_TK[31]:B 
*.PININFO WL_TK[32]:B WL_TK[33]:B WL_TK[34]:B WL_TK[35]:B WL_TK[36]:B 
*.PININFO WL_TK[37]:B WL_TK[38]:B WL_TK[39]:B WL_TK[40]:B WL_TK[41]:B 
*.PININFO WL_TK[42]:B WL_TK[43]:B WL_TK[44]:B WL_TK[45]:B WL_TK[46]:B 
*.PININFO WL_TK[47]:B WL_TK[48]:B WL_TK[49]:B WL_TK[50]:B WL_TK[51]:B 
*.PININFO WL_TK[52]:B WL_TK[53]:B WL_TK[54]:B WL_TK[55]:B WL_TK[56]:B 
*.PININFO WL_TK[57]:B WL_TK[58]:B WL_TK[59]:B WL_TK[60]:B WL_TK[61]:B 
*.PININFO WL_TK[62]:B WL_TK[63]:B WL_TK[64]:B WL_TK[65]:B WL_TK[66]:B 
*.PININFO WL_TK[67]:B WL_TK[68]:B WL_TK[69]:B WL_TK[70]:B WL_TK[71]:B 
*.PININFO WL_TK[72]:B WL_TK[73]:B WL_TK[74]:B WL_TK[75]:B WL_TK[76]:B 
*.PININFO WL_TK[77]:B WL_TK[78]:B WL_TK[79]:B WL_TK[80]:B WL_TK[81]:B 
*.PININFO WL_TK[82]:B WL_TK[83]:B WL_TK[84]:B WL_TK[85]:B WL_TK[86]:B 
*.PININFO WL_TK[87]:B WL_TK[88]:B WL_TK[89]:B WL_TK[90]:B WL_TK[91]:B 
*.PININFO WL_TK[92]:B WL_TK[93]:B WL_TK[94]:B WL_TK[95]:B WL_TK[96]:B 
*.PININFO WL_TK[97]:B WL_TK[98]:B WL_TK[99]:B WL_TK[100]:B WL_TK[101]:B 
*.PININFO WL_TK[102]:B WL_TK[103]:B WL_TK[104]:B WL_TK[105]:B WL_TK[106]:B 
*.PININFO WL_TK[107]:B WL_TK[108]:B WL_TK[109]:B WL_TK[110]:B WL_TK[111]:B 
*.PININFO WL_TK[112]:B WL_TK[113]:B WL_TK[114]:B WL_TK[115]:B WL_TK[116]:B 
*.PININFO WL_TK[117]:B WL_TK[118]:B WL_TK[119]:B WL_TK[120]:B WL_TK[121]:B 
*.PININFO WL_TK[122]:B WL_TK[123]:B WL_TK[124]:B WL_TK[125]:B WL_TK[126]:B 
*.PININFO WL_TK[127]:B WL_TK[128]:B WL_TK[129]:B WL_TK[130]:B WL_TK[131]:B 
*.PININFO WL_TK[132]:B WL_TK[133]:B WL_TK[134]:B WL_TK[135]:B WL_TK[136]:B 
*.PININFO WL_TK[137]:B WL_TK[138]:B WL_TK[139]:B WL_TK[140]:B WL_TK[141]:B 
*.PININFO WL_TK[142]:B WL_TK[143]:B WL_TK[144]:B WL_TK[145]:B WL_TK[146]:B 
*.PININFO WL_TK[147]:B WL_TK[148]:B WL_TK[149]:B WL_TK[150]:B WL_TK[151]:B 
*.PININFO WL_TK[152]:B WL_TK[153]:B WL_TK[154]:B WL_TK[155]:B WL_TK[156]:B 
*.PININFO WL_TK[157]:B WL_TK[158]:B WL_TK[159]:B WL_TK[160]:B WL_TK[161]:B 
*.PININFO WL_TK[162]:B WL_TK[163]:B WL_TK[164]:B WL_TK[165]:B WL_TK[166]:B 
*.PININFO WL_TK[167]:B WL_TK[168]:B WL_TK[169]:B WL_TK[170]:B WL_TK[171]:B 
*.PININFO WL_TK[172]:B WL_TK[173]:B WL_TK[174]:B WL_TK[175]:B WL_TK[176]:B 
*.PININFO WL_TK[177]:B WL_TK[178]:B WL_TK[179]:B WL_TK[180]:B WL_TK[181]:B 
*.PININFO WL_TK[182]:B WL_TK[183]:B WL_TK[184]:B WL_TK[185]:B WL_TK[186]:B 
*.PININFO WL_TK[187]:B WL_TK[188]:B WL_TK[189]:B WL_TK[190]:B WL_TK[191]:B 
*.PININFO WL_TK[192]:B WL_TK[193]:B WL_TK[194]:B WL_TK[195]:B WL_TK[196]:B 
*.PININFO WL_TK[197]:B WL_TK[198]:B WL_TK[199]:B WL_TK[200]:B WL_TK[201]:B 
*.PININFO WL_TK[202]:B WL_TK[203]:B WL_TK[204]:B WL_TK[205]:B WL_TK[206]:B 
*.PININFO WL_TK[207]:B WL_TK[208]:B WL_TK[209]:B WL_TK[210]:B WL_TK[211]:B 
*.PININFO WL_TK[212]:B WL_TK[213]:B WL_TK[214]:B WL_TK[215]:B WL_TK[216]:B 
*.PININFO WL_TK[217]:B WL_TK[218]:B WL_TK[219]:B WL_TK[220]:B WL_TK[221]:B 
*.PININFO WL_TK[222]:B WL_TK[223]:B WL_TK[224]:B WL_TK[225]:B WL_TK[226]:B 
*.PININFO WL_TK[227]:B WL_TK[228]:B WL_TK[229]:B WL_TK[230]:B WL_TK[231]:B 
*.PININFO WL_TK[232]:B WL_TK[233]:B WL_TK[234]:B WL_TK[235]:B WL_TK[236]:B 
*.PININFO WL_TK[237]:B WL_TK[238]:B WL_TK[239]:B WL_TK[240]:B WL_TK[241]:B 
*.PININFO WL_TK[242]:B WL_TK[243]:B WL_TK[244]:B WL_TK[245]:B WL_TK[246]:B 
*.PININFO WL_TK[247]:B WL_TK[248]:B WL_TK[249]:B WL_TK[250]:B WL_TK[251]:B 
*.PININFO WL_TK[252]:B WL_TK[253]:B WL_TK[254]:B WL_TK[255]:B WL_TK[256]:B 
*.PININFO WL_TK[257]:B WL_TK[258]:B WL_TK[259]:B WL_TK[260]:B WL_TK[261]:B 
*.PININFO WL_TK[262]:B WL_TK[263]:B WL_TK[264]:B WL_TK[265]:B WL_TK[266]:B 
*.PININFO WL_TK[267]:B WL_TK[268]:B WL_TK[269]:B WL_TK[270]:B WL_TK[271]:B 
*.PININFO WL_TK[272]:B WL_TK[273]:B WL_TK[274]:B WL_TK[275]:B WL_TK[276]:B 
*.PININFO WL_TK[277]:B WL_TK[278]:B WL_TK[279]:B WL_TK[280]:B WL_TK[281]:B 
*.PININFO WL_TK[282]:B WL_TK[283]:B WL_TK[284]:B WL_TK[285]:B WL_TK[286]:B 
*.PININFO WL_TK[287]:B WL_TK[288]:B WL_TK[289]:B WL_TK[290]:B WL_TK[291]:B 
*.PININFO WL_TK[292]:B WL_TK[293]:B WL_TK[294]:B WL_TK[295]:B WL_TK[296]:B 
*.PININFO WL_TK[297]:B WL_TK[298]:B WL_TK[299]:B WL_TK[300]:B WL_TK[301]:B 
*.PININFO WL_TK[302]:B WL_TK[303]:B WL_TK[304]:B WL_TK[305]:B WL_TK[306]:B 
*.PININFO WL_TK[307]:B WL_TK[308]:B WL_TK[309]:B WL_TK[310]:B WL_TK[311]:B 
*.PININFO WL_TK[312]:B WL_TK[313]:B WL_TK[314]:B WL_TK[315]:B WL_TK[316]:B 
*.PININFO WL_TK[317]:B WL_TK[318]:B WL_TK[319]:B WL_TK[320]:B WL_TK[321]:B 
*.PININFO WL_TK[322]:B WL_TK[323]:B WL_TK[324]:B WL_TK[325]:B WL_TK[326]:B 
*.PININFO WL_TK[327]:B WL_TK[328]:B WL_TK[329]:B WL_TK[330]:B WL_TK[331]:B 
*.PININFO WL_TK[332]:B WL_TK[333]:B WL_TK[334]:B WL_TK[335]:B WL_TK[336]:B 
*.PININFO WL_TK[337]:B WL_TK[338]:B WL_TK[339]:B WL_TK[340]:B WL_TK[341]:B 
*.PININFO WL_TK[342]:B WL_TK[343]:B WL_TK[344]:B WL_TK[345]:B WL_TK[346]:B 
*.PININFO WL_TK[347]:B WL_TK[348]:B WL_TK[349]:B WL_TK[350]:B WL_TK[351]:B 
*.PININFO WL_TK[352]:B WL_TK[353]:B WL_TK[354]:B WL_TK[355]:B WL_TK[356]:B 
*.PININFO WL_TK[357]:B WL_TK[358]:B WL_TK[359]:B WL_TK[360]:B WL_TK[361]:B 
*.PININFO WL_TK[362]:B WL_TK[363]:B WL_TK[364]:B WL_TK[365]:B WL_TK[366]:B 
*.PININFO WL_TK[367]:B WL_TK[368]:B WL_TK[369]:B WL_TK[370]:B WL_TK[371]:B 
*.PININFO WL_TK[372]:B WL_TK[373]:B WL_TK[374]:B WL_TK[375]:B WL_TK[376]:B 
*.PININFO WL_TK[377]:B WL_TK[378]:B WL_TK[379]:B WL_TK[380]:B WL_TK[381]:B 
*.PININFO WL_TK[382]:B WL_TK[383]:B WL_TK[384]:B WL_TK[385]:B WL_TK[386]:B 
*.PININFO WL_TK[387]:B WL_TK[388]:B WL_TK[389]:B WL_TK[390]:B WL_TK[391]:B 
*.PININFO WL_TK[392]:B WL_TK[393]:B WL_TK[394]:B WL_TK[395]:B WL_TK[396]:B 
*.PININFO WL_TK[397]:B WL_TK[398]:B WL_TK[399]:B WL_TK[400]:B WL_TK[401]:B 
*.PININFO WL_TK[402]:B WL_TK[403]:B WL_TK[404]:B WL_TK[405]:B WL_TK[406]:B 
*.PININFO WL_TK[407]:B WL_TK[408]:B WL_TK[409]:B WL_TK[410]:B WL_TK[411]:B 
*.PININFO WL_TK[412]:B WL_TK[413]:B WL_TK[414]:B WL_TK[415]:B WL_TK[416]:B 
*.PININFO WL_TK[417]:B WL_TK[418]:B WL_TK[419]:B WL_TK[420]:B WL_TK[421]:B 
*.PININFO WL_TK[422]:B WL_TK[423]:B WL_TK[424]:B WL_TK[425]:B WL_TK[426]:B 
*.PININFO WL_TK[427]:B WL_TK[428]:B WL_TK[429]:B WL_TK[430]:B WL_TK[431]:B 
*.PININFO WL_TK[432]:B WL_TK[433]:B WL_TK[434]:B WL_TK[435]:B WL_TK[436]:B 
*.PININFO WL_TK[437]:B WL_TK[438]:B WL_TK[439]:B WL_TK[440]:B WL_TK[441]:B 
*.PININFO WL_TK[442]:B WL_TK[443]:B WL_TK[444]:B WL_TK[445]:B WL_TK[446]:B 
*.PININFO WL_TK[447]:B WL_TK[448]:B WL_TK[449]:B WL_TK[450]:B WL_TK[451]:B 
*.PININFO WL_TK[452]:B WL_TK[453]:B WL_TK[454]:B WL_TK[455]:B WL_TK[456]:B 
*.PININFO WL_TK[457]:B WL_TK[458]:B WL_TK[459]:B WL_TK[460]:B WL_TK[461]:B 
*.PININFO WL_TK[462]:B WL_TK[463]:B WL_TK[464]:B WL_TK[465]:B WL_TK[466]:B 
*.PININFO WL_TK[467]:B WL_TK[468]:B WL_TK[469]:B WL_TK[470]:B WL_TK[471]:B 
*.PININFO WL_TK[472]:B WL_TK[473]:B WL_TK[474]:B WL_TK[475]:B WL_TK[476]:B 
*.PININFO WL_TK[477]:B WL_TK[478]:B WL_TK[479]:B WL_TK[480]:B WL_TK[481]:B 
*.PININFO WL_TK[482]:B WL_TK[483]:B WL_TK[484]:B WL_TK[485]:B WL_TK[486]:B 
*.PININFO WL_TK[487]:B WL_TK[488]:B WL_TK[489]:B WL_TK[490]:B WL_TK[491]:B 
*.PININFO WL_TK[492]:B WL_TK[493]:B WL_TK[494]:B WL_TK[495]:B WL_TK[496]:B 
*.PININFO WL_TK[497]:B WL_TK[498]:B WL_TK[499]:B WL_TK[500]:B WL_TK[501]:B 
*.PININFO WL_TK[502]:B WL_TK[503]:B WL_TK[504]:B WL_TK[505]:B WL_TK[506]:B 
*.PININFO WL_TK[507]:B WL_TK[508]:B WL_TK[509]:B WL_TK[510]:B WL_TK[511]:B 
*.PININFO TIEH:B TIEL:B
XTRKNORX64_DUMY6 BL_TK VDDI VSSI WL[256] WL[257] WL[258] WL[259] WL[260] 
+ WL[261] WL[262] WL[263] WL[264] WL[265] WL[266] WL[267] WL[268] WL[269] 
+ WL[270] WL[271] WL[272] WL[273] WL[274] WL[275] WL[276] WL[277] WL[278] 
+ WL[279] WL[280] WL[281] WL[282] WL[283] WL[284] WL[285] WL[286] WL[287] 
+ WL[288] WL[289] WL[290] WL[291] WL[292] WL[293] WL[294] WL[295] WL[296] 
+ WL[297] WL[298] WL[299] WL[300] WL[301] WL[302] WL[303] WL[304] WL[305] 
+ WL[306] WL[307] WL[308] WL[309] WL[310] WL[311] WL[312] WL[313] WL[314] 
+ WL[315] WL[316] WL[317] WL[318] WL[319] WL_TK[256] WL_TK[257] WL_TK[258] 
+ WL_TK[259] WL_TK[260] WL_TK[261] WL_TK[262] WL_TK[263] WL_TK[264] WL_TK[265] 
+ WL_TK[266] WL_TK[267] WL_TK[268] WL_TK[269] WL_TK[270] WL_TK[271] WL_TK[272] 
+ WL_TK[273] WL_TK[274] WL_TK[275] WL_TK[276] WL_TK[277] WL_TK[278] WL_TK[279] 
+ WL_TK[280] WL_TK[281] WL_TK[282] WL_TK[283] WL_TK[284] WL_TK[285] WL_TK[286] 
+ WL_TK[287] WL_TK[288] WL_TK[289] WL_TK[290] WL_TK[291] WL_TK[292] WL_TK[293] 
+ WL_TK[294] WL_TK[295] WL_TK[296] WL_TK[297] WL_TK[298] WL_TK[299] WL_TK[300] 
+ WL_TK[301] WL_TK[302] WL_TK[303] WL_TK[304] WL_TK[305] WL_TK[306] WL_TK[307] 
+ WL_TK[308] WL_TK[309] WL_TK[310] WL_TK[311] WL_TK[312] WL_TK[313] WL_TK[314] 
+ WL_TK[315] WL_TK[316] WL_TK[317] WL_TK[318] WL_TK[319] NET49[0] NET49[1] 
+ NET49[2] NET49[3] NET49[4] NET49[5] NET49[6] NET49[7] NET49[8] NET49[9] 
+ NET49[10] NET49[11] NET49[12] NET49[13] NET49[14] NET49[15] NET49[16] 
+ NET49[17] NET49[18] NET49[19] NET49[20] NET49[21] NET49[22] NET49[23] 
+ NET49[24] NET49[25] NET49[26] NET49[27] NET49[28] NET49[29] NET49[30] 
+ NET49[31] NET48 NET47 NET46[0] NET46[1] NET46[2] NET46[3] NET46[4] NET46[5] 
+ NET46[6] NET46[7] NET46[8] NET46[9] NET46[10] NET46[11] NET46[12] NET46[13] 
+ NET46[14] NET46[15] NET46[16] NET46[17] NET46[18] NET46[19] NET46[20] 
+ NET46[21] NET46[22] NET46[23] NET46[24] NET46[25] NET46[26] NET46[27] 
+ NET46[28] NET46[29] NET46[30] NET46[31] TIEH S1AHSF400W40_TRKNORX64_CHAR
XTRKNORX64_DUMY4 BL_TK VDDI VSSI WL[128] WL[129] WL[130] WL[131] WL[132] 
+ WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] WL[140] WL[141] 
+ WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] WL[149] WL[150] 
+ WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] WL[158] WL[159] 
+ WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] WL[167] WL[168] 
+ WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] WL[176] WL[177] 
+ WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] WL[185] WL[186] 
+ WL[187] WL[188] WL[189] WL[190] WL[191] WL_TK[128] WL_TK[129] WL_TK[130] 
+ WL_TK[131] WL_TK[132] WL_TK[133] WL_TK[134] WL_TK[135] WL_TK[136] WL_TK[137] 
+ WL_TK[138] WL_TK[139] WL_TK[140] WL_TK[141] WL_TK[142] WL_TK[143] WL_TK[144] 
+ WL_TK[145] WL_TK[146] WL_TK[147] WL_TK[148] WL_TK[149] WL_TK[150] WL_TK[151] 
+ WL_TK[152] WL_TK[153] WL_TK[154] WL_TK[155] WL_TK[156] WL_TK[157] WL_TK[158] 
+ WL_TK[159] WL_TK[160] WL_TK[161] WL_TK[162] WL_TK[163] WL_TK[164] WL_TK[165] 
+ WL_TK[166] WL_TK[167] WL_TK[168] WL_TK[169] WL_TK[170] WL_TK[171] WL_TK[172] 
+ WL_TK[173] WL_TK[174] WL_TK[175] WL_TK[176] WL_TK[177] WL_TK[178] WL_TK[179] 
+ WL_TK[180] WL_TK[181] WL_TK[182] WL_TK[183] WL_TK[184] WL_TK[185] WL_TK[186] 
+ WL_TK[187] WL_TK[188] WL_TK[189] WL_TK[190] WL_TK[191] NET59[0] NET59[1] 
+ NET59[2] NET59[3] NET59[4] NET59[5] NET59[6] NET59[7] NET59[8] NET59[9] 
+ NET59[10] NET59[11] NET59[12] NET59[13] NET59[14] NET59[15] NET59[16] 
+ NET59[17] NET59[18] NET59[19] NET59[20] NET59[21] NET59[22] NET59[23] 
+ NET59[24] NET59[25] NET59[26] NET59[27] NET59[28] NET59[29] NET59[30] 
+ NET59[31] NET58 NET57 NET56[0] NET56[1] NET56[2] NET56[3] NET56[4] NET56[5] 
+ NET56[6] NET56[7] NET56[8] NET56[9] NET56[10] NET56[11] NET56[12] NET56[13] 
+ NET56[14] NET56[15] NET56[16] NET56[17] NET56[18] NET56[19] NET56[20] 
+ NET56[21] NET56[22] NET56[23] NET56[24] NET56[25] NET56[26] NET56[27] 
+ NET56[28] NET56[29] NET56[30] NET56[31] TIEH S1AHSF400W40_TRKNORX64_CHAR
XTRKNORX64_DUMY7 BL_TK VDDI VSSI WL[320] WL[321] WL[322] WL[323] WL[324] 
+ WL[325] WL[326] WL[327] WL[328] WL[329] WL[330] WL[331] WL[332] WL[333] 
+ WL[334] WL[335] WL[336] WL[337] WL[338] WL[339] WL[340] WL[341] WL[342] 
+ WL[343] WL[344] WL[345] WL[346] WL[347] WL[348] WL[349] WL[350] WL[351] 
+ WL[352] WL[353] WL[354] WL[355] WL[356] WL[357] WL[358] WL[359] WL[360] 
+ WL[361] WL[362] WL[363] WL[364] WL[365] WL[366] WL[367] WL[368] WL[369] 
+ WL[370] WL[371] WL[372] WL[373] WL[374] WL[375] WL[376] WL[377] WL[378] 
+ WL[379] WL[380] WL[381] WL[382] WL[383] WL_TK[320] WL_TK[321] WL_TK[322] 
+ WL_TK[323] WL_TK[324] WL_TK[325] WL_TK[326] WL_TK[327] WL_TK[328] WL_TK[329] 
+ WL_TK[330] WL_TK[331] WL_TK[332] WL_TK[333] WL_TK[334] WL_TK[335] WL_TK[336] 
+ WL_TK[337] WL_TK[338] WL_TK[339] WL_TK[340] WL_TK[341] WL_TK[342] WL_TK[343] 
+ WL_TK[344] WL_TK[345] WL_TK[346] WL_TK[347] WL_TK[348] WL_TK[349] WL_TK[350] 
+ WL_TK[351] WL_TK[352] WL_TK[353] WL_TK[354] WL_TK[355] WL_TK[356] WL_TK[357] 
+ WL_TK[358] WL_TK[359] WL_TK[360] WL_TK[361] WL_TK[362] WL_TK[363] WL_TK[364] 
+ WL_TK[365] WL_TK[366] WL_TK[367] WL_TK[368] WL_TK[369] WL_TK[370] WL_TK[371] 
+ WL_TK[372] WL_TK[373] WL_TK[374] WL_TK[375] WL_TK[376] WL_TK[377] WL_TK[378] 
+ WL_TK[379] WL_TK[380] WL_TK[381] WL_TK[382] WL_TK[383] NET39[0] NET39[1] 
+ NET39[2] NET39[3] NET39[4] NET39[5] NET39[6] NET39[7] NET39[8] NET39[9] 
+ NET39[10] NET39[11] NET39[12] NET39[13] NET39[14] NET39[15] NET39[16] 
+ NET39[17] NET39[18] NET39[19] NET39[20] NET39[21] NET39[22] NET39[23] 
+ NET39[24] NET39[25] NET39[26] NET39[27] NET39[28] NET39[29] NET39[30] 
+ NET39[31] NET38 NET37 NET36[0] NET36[1] NET36[2] NET36[3] NET36[4] NET36[5] 
+ NET36[6] NET36[7] NET36[8] NET36[9] NET36[10] NET36[11] NET36[12] NET36[13] 
+ NET36[14] NET36[15] NET36[16] NET36[17] NET36[18] NET36[19] NET36[20] 
+ NET36[21] NET36[22] NET36[23] NET36[24] NET36[25] NET36[26] NET36[27] 
+ NET36[28] NET36[29] NET36[30] NET36[31] TIEH S1AHSF400W40_TRKNORX64_CHAR
XTRKNORX64_DUMY3 BL_TK VDDI VSSI WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] 
+ WL[70] WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] 
+ WL[81] WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] 
+ WL[92] WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] 
+ WL[102] WL[103] WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] 
+ WL[111] WL[112] WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] 
+ WL[120] WL[121] WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL_TK[64] 
+ WL_TK[65] WL_TK[66] WL_TK[67] WL_TK[68] WL_TK[69] WL_TK[70] WL_TK[71] 
+ WL_TK[72] WL_TK[73] WL_TK[74] WL_TK[75] WL_TK[76] WL_TK[77] WL_TK[78] 
+ WL_TK[79] WL_TK[80] WL_TK[81] WL_TK[82] WL_TK[83] WL_TK[84] WL_TK[85] 
+ WL_TK[86] WL_TK[87] WL_TK[88] WL_TK[89] WL_TK[90] WL_TK[91] WL_TK[92] 
+ WL_TK[93] WL_TK[94] WL_TK[95] WL_TK[96] WL_TK[97] WL_TK[98] WL_TK[99] 
+ WL_TK[100] WL_TK[101] WL_TK[102] WL_TK[103] WL_TK[104] WL_TK[105] WL_TK[106] 
+ WL_TK[107] WL_TK[108] WL_TK[109] WL_TK[110] WL_TK[111] WL_TK[112] WL_TK[113] 
+ WL_TK[114] WL_TK[115] WL_TK[116] WL_TK[117] WL_TK[118] WL_TK[119] WL_TK[120] 
+ WL_TK[121] WL_TK[122] WL_TK[123] WL_TK[124] WL_TK[125] WL_TK[126] WL_TK[127] 
+ NET69[0] NET69[1] NET69[2] NET69[3] NET69[4] NET69[5] NET69[6] NET69[7] 
+ NET69[8] NET69[9] NET69[10] NET69[11] NET69[12] NET69[13] NET69[14] 
+ NET69[15] NET69[16] NET69[17] NET69[18] NET69[19] NET69[20] NET69[21] 
+ NET69[22] NET69[23] NET69[24] NET69[25] NET69[26] NET69[27] NET69[28] 
+ NET69[29] NET69[30] NET69[31] NET68 NET67 NET66[0] NET66[1] NET66[2] 
+ NET66[3] NET66[4] NET66[5] NET66[6] NET66[7] NET66[8] NET66[9] NET66[10] 
+ NET66[11] NET66[12] NET66[13] NET66[14] NET66[15] NET66[16] NET66[17] 
+ NET66[18] NET66[19] NET66[20] NET66[21] NET66[22] NET66[23] NET66[24] 
+ NET66[25] NET66[26] NET66[27] NET66[28] NET66[29] NET66[30] NET66[31] TIEH 
+ S1AHSF400W40_TRKNORX64_CHAR
XTRKNORX64_DYMY5 BL_TK VDDI VSSI WL[192] WL[193] WL[194] WL[195] WL[196] 
+ WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] WL[203] WL[204] WL[205] 
+ WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] WL[212] WL[213] WL[214] 
+ WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] WL[221] WL[222] WL[223] 
+ WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] WL[230] WL[231] WL[232] 
+ WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] WL[239] WL[240] WL[241] 
+ WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] WL[248] WL[249] WL[250] 
+ WL[251] WL[252] WL[253] WL[254] WL[255] WL_TK[192] WL_TK[193] WL_TK[194] 
+ WL_TK[195] WL_TK[196] WL_TK[197] WL_TK[198] WL_TK[199] WL_TK[200] WL_TK[201] 
+ WL_TK[202] WL_TK[203] WL_TK[204] WL_TK[205] WL_TK[206] WL_TK[207] WL_TK[208] 
+ WL_TK[209] WL_TK[210] WL_TK[211] WL_TK[212] WL_TK[213] WL_TK[214] WL_TK[215] 
+ WL_TK[216] WL_TK[217] WL_TK[218] WL_TK[219] WL_TK[220] WL_TK[221] WL_TK[222] 
+ WL_TK[223] WL_TK[224] WL_TK[225] WL_TK[226] WL_TK[227] WL_TK[228] WL_TK[229] 
+ WL_TK[230] WL_TK[231] WL_TK[232] WL_TK[233] WL_TK[234] WL_TK[235] WL_TK[236] 
+ WL_TK[237] WL_TK[238] WL_TK[239] WL_TK[240] WL_TK[241] WL_TK[242] WL_TK[243] 
+ WL_TK[244] WL_TK[245] WL_TK[246] WL_TK[247] WL_TK[248] WL_TK[249] WL_TK[250] 
+ WL_TK[251] WL_TK[252] WL_TK[253] WL_TK[254] WL_TK[255] NET79[0] NET79[1] 
+ NET79[2] NET79[3] NET79[4] NET79[5] NET79[6] NET79[7] NET79[8] NET79[9] 
+ NET79[10] NET79[11] NET79[12] NET79[13] NET79[14] NET79[15] NET79[16] 
+ NET79[17] NET79[18] NET79[19] NET79[20] NET79[21] NET79[22] NET79[23] 
+ NET79[24] NET79[25] NET79[26] NET79[27] NET79[28] NET79[29] NET79[30] 
+ NET79[31] NET78 NET77 NET76[0] NET76[1] NET76[2] NET76[3] NET76[4] NET76[5] 
+ NET76[6] NET76[7] NET76[8] NET76[9] NET76[10] NET76[11] NET76[12] NET76[13] 
+ NET76[14] NET76[15] NET76[16] NET76[17] NET76[18] NET76[19] NET76[20] 
+ NET76[21] NET76[22] NET76[23] NET76[24] NET76[25] NET76[26] NET76[27] 
+ NET76[28] NET76[29] NET76[30] NET76[31] TIEH S1AHSF400W40_TRKNORX64_CHAR
XTRKNORX16_DUMY0 BL_TK VDDI VSSI WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] 
+ WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] 
+ WL_TK[16] WL_TK[17] WL_TK[18] WL_TK[19] WL_TK[20] WL_TK[21] WL_TK[22] 
+ WL_TK[23] WL_TK[24] WL_TK[25] WL_TK[26] WL_TK[27] WL_TK[28] WL_TK[29] 
+ WL_TK[30] WL_TK[31] NET89[0] NET89[1] NET89[2] NET89[3] NET89[4] NET89[5] 
+ NET89[6] NET89[7] NET88 NET108 NET86[0] NET86[1] NET86[2] NET86[3] NET86[4] 
+ NET86[5] NET86[6] NET86[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
XTRKNORX16_DUMY1 BL_TK VDDI VSSI WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] 
+ WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] 
+ WL_TK[32] WL_TK[33] WL_TK[34] WL_TK[35] WL_TK[36] WL_TK[37] WL_TK[38] 
+ WL_TK[39] WL_TK[40] WL_TK[41] WL_TK[42] WL_TK[43] WL_TK[44] WL_TK[45] 
+ WL_TK[46] WL_TK[47] NET99[0] NET99[1] NET99[2] NET99[3] NET99[4] NET99[5] 
+ NET99[6] NET99[7] NET98 NET88 NET96[0] NET96[1] NET96[2] NET96[3] NET96[4] 
+ NET96[5] NET96[6] NET96[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
XTRKNORX16_BCELL BL_TK VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] 
+ WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL_TK[0] 
+ WL_TK[1] WL_TK[2] WL_TK[3] WL_TK[4] WL_TK[5] WL_TK[6] WL_TK[7] WL_TK[8] 
+ WL_TK[9] WL_TK[10] WL_TK[11] WL_TK[12] WL_TK[13] WL_TK[14] WL_TK[15] 
+ NET109[0] NET109[1] NET109[2] NET109[3] NET109[4] NET109[5] NET109[6] 
+ NET109[7] NET108 NET107 NET106[0] NET106[1] NET106[2] NET106[3] NET106[4] 
+ NET106[5] NET106[6] NET106[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
XTRKNORX16_DUMY2 BL_TK VDDI VSSI WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] 
+ WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] 
+ WL_TK[48] WL_TK[49] WL_TK[50] WL_TK[51] WL_TK[52] WL_TK[53] WL_TK[54] 
+ WL_TK[55] WL_TK[56] WL_TK[57] WL_TK[58] WL_TK[59] WL_TK[60] WL_TK[61] 
+ WL_TK[62] WL_TK[63] NET119[0] NET119[1] NET119[2] NET119[3] NET119[4] 
+ NET119[5] NET119[6] NET119[7] NET118 NET98 NET116[0] NET116[1] NET116[2] 
+ NET116[3] NET116[4] NET116[5] NET116[6] NET116[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    TKBL_S512_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TKBL_S512_CHAR BL_TK VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] WL_TK[0] WL_TK[1] WL_TK[2] WL_TK[3] WL_TK[4] 
+ WL_TK[5] WL_TK[6] WL_TK[7] WL_TK[8] WL_TK[9] WL_TK[10] WL_TK[11] WL_TK[12] 
+ WL_TK[13] WL_TK[14] WL_TK[15] WL_TK[16] WL_TK[17] WL_TK[18] WL_TK[19] 
+ WL_TK[20] WL_TK[21] WL_TK[22] WL_TK[23] WL_TK[24] WL_TK[25] WL_TK[26] 
+ WL_TK[27] WL_TK[28] WL_TK[29] WL_TK[30] WL_TK[31] WL_TK[32] WL_TK[33] 
+ WL_TK[34] WL_TK[35] WL_TK[36] WL_TK[37] WL_TK[38] WL_TK[39] WL_TK[40] 
+ WL_TK[41] WL_TK[42] WL_TK[43] WL_TK[44] WL_TK[45] WL_TK[46] WL_TK[47] 
+ WL_TK[48] WL_TK[49] WL_TK[50] WL_TK[51] WL_TK[52] WL_TK[53] WL_TK[54] 
+ WL_TK[55] WL_TK[56] WL_TK[57] WL_TK[58] WL_TK[59] WL_TK[60] WL_TK[61] 
+ WL_TK[62] WL_TK[63] WL_TK[64] WL_TK[65] WL_TK[66] WL_TK[67] WL_TK[68] 
+ WL_TK[69] WL_TK[70] WL_TK[71] WL_TK[72] WL_TK[73] WL_TK[74] WL_TK[75] 
+ WL_TK[76] WL_TK[77] WL_TK[78] WL_TK[79] WL_TK[80] WL_TK[81] WL_TK[82] 
+ WL_TK[83] WL_TK[84] WL_TK[85] WL_TK[86] WL_TK[87] WL_TK[88] WL_TK[89] 
+ WL_TK[90] WL_TK[91] WL_TK[92] WL_TK[93] WL_TK[94] WL_TK[95] WL_TK[96] 
+ WL_TK[97] WL_TK[98] WL_TK[99] WL_TK[100] WL_TK[101] WL_TK[102] WL_TK[103] 
+ WL_TK[104] WL_TK[105] WL_TK[106] WL_TK[107] WL_TK[108] WL_TK[109] WL_TK[110] 
+ WL_TK[111] WL_TK[112] WL_TK[113] WL_TK[114] WL_TK[115] WL_TK[116] WL_TK[117] 
+ WL_TK[118] WL_TK[119] WL_TK[120] WL_TK[121] WL_TK[122] WL_TK[123] WL_TK[124] 
+ WL_TK[125] WL_TK[126] WL_TK[127] WL_TK[128] WL_TK[129] WL_TK[130] WL_TK[131] 
+ WL_TK[132] WL_TK[133] WL_TK[134] WL_TK[135] WL_TK[136] WL_TK[137] WL_TK[138] 
+ WL_TK[139] WL_TK[140] WL_TK[141] WL_TK[142] WL_TK[143] WL_TK[144] WL_TK[145] 
+ WL_TK[146] WL_TK[147] WL_TK[148] WL_TK[149] WL_TK[150] WL_TK[151] WL_TK[152] 
+ WL_TK[153] WL_TK[154] WL_TK[155] WL_TK[156] WL_TK[157] WL_TK[158] WL_TK[159] 
+ WL_TK[160] WL_TK[161] WL_TK[162] WL_TK[163] WL_TK[164] WL_TK[165] WL_TK[166] 
+ WL_TK[167] WL_TK[168] WL_TK[169] WL_TK[170] WL_TK[171] WL_TK[172] WL_TK[173] 
+ WL_TK[174] WL_TK[175] WL_TK[176] WL_TK[177] WL_TK[178] WL_TK[179] WL_TK[180] 
+ WL_TK[181] WL_TK[182] WL_TK[183] WL_TK[184] WL_TK[185] WL_TK[186] WL_TK[187] 
+ WL_TK[188] WL_TK[189] WL_TK[190] WL_TK[191] WL_TK[192] WL_TK[193] WL_TK[194] 
+ WL_TK[195] WL_TK[196] WL_TK[197] WL_TK[198] WL_TK[199] WL_TK[200] WL_TK[201] 
+ WL_TK[202] WL_TK[203] WL_TK[204] WL_TK[205] WL_TK[206] WL_TK[207] WL_TK[208] 
+ WL_TK[209] WL_TK[210] WL_TK[211] WL_TK[212] WL_TK[213] WL_TK[214] WL_TK[215] 
+ WL_TK[216] WL_TK[217] WL_TK[218] WL_TK[219] WL_TK[220] WL_TK[221] WL_TK[222] 
+ WL_TK[223] WL_TK[224] WL_TK[225] WL_TK[226] WL_TK[227] WL_TK[228] WL_TK[229] 
+ WL_TK[230] WL_TK[231] WL_TK[232] WL_TK[233] WL_TK[234] WL_TK[235] WL_TK[236] 
+ WL_TK[237] WL_TK[238] WL_TK[239] WL_TK[240] WL_TK[241] WL_TK[242] WL_TK[243] 
+ WL_TK[244] WL_TK[245] WL_TK[246] WL_TK[247] WL_TK[248] WL_TK[249] WL_TK[250] 
+ WL_TK[251] WL_TK[252] WL_TK[253] WL_TK[254] WL_TK[255] WL_TK[256] WL_TK[257] 
+ WL_TK[258] WL_TK[259] WL_TK[260] WL_TK[261] WL_TK[262] WL_TK[263] WL_TK[264] 
+ WL_TK[265] WL_TK[266] WL_TK[267] WL_TK[268] WL_TK[269] WL_TK[270] WL_TK[271] 
+ WL_TK[272] WL_TK[273] WL_TK[274] WL_TK[275] WL_TK[276] WL_TK[277] WL_TK[278] 
+ WL_TK[279] WL_TK[280] WL_TK[281] WL_TK[282] WL_TK[283] WL_TK[284] WL_TK[285] 
+ WL_TK[286] WL_TK[287] WL_TK[288] WL_TK[289] WL_TK[290] WL_TK[291] WL_TK[292] 
+ WL_TK[293] WL_TK[294] WL_TK[295] WL_TK[296] WL_TK[297] WL_TK[298] WL_TK[299] 
+ WL_TK[300] WL_TK[301] WL_TK[302] WL_TK[303] WL_TK[304] WL_TK[305] WL_TK[306] 
+ WL_TK[307] WL_TK[308] WL_TK[309] WL_TK[310] WL_TK[311] WL_TK[312] WL_TK[313] 
+ WL_TK[314] WL_TK[315] WL_TK[316] WL_TK[317] WL_TK[318] WL_TK[319] WL_TK[320] 
+ WL_TK[321] WL_TK[322] WL_TK[323] WL_TK[324] WL_TK[325] WL_TK[326] WL_TK[327] 
+ WL_TK[328] WL_TK[329] WL_TK[330] WL_TK[331] WL_TK[332] WL_TK[333] WL_TK[334] 
+ WL_TK[335] WL_TK[336] WL_TK[337] WL_TK[338] WL_TK[339] WL_TK[340] WL_TK[341] 
+ WL_TK[342] WL_TK[343] WL_TK[344] WL_TK[345] WL_TK[346] WL_TK[347] WL_TK[348] 
+ WL_TK[349] WL_TK[350] WL_TK[351] WL_TK[352] WL_TK[353] WL_TK[354] WL_TK[355] 
+ WL_TK[356] WL_TK[357] WL_TK[358] WL_TK[359] WL_TK[360] WL_TK[361] WL_TK[362] 
+ WL_TK[363] WL_TK[364] WL_TK[365] WL_TK[366] WL_TK[367] WL_TK[368] WL_TK[369] 
+ WL_TK[370] WL_TK[371] WL_TK[372] WL_TK[373] WL_TK[374] WL_TK[375] WL_TK[376] 
+ WL_TK[377] WL_TK[378] WL_TK[379] WL_TK[380] WL_TK[381] WL_TK[382] WL_TK[383] 
+ WL_TK[384] WL_TK[385] WL_TK[386] WL_TK[387] WL_TK[388] WL_TK[389] WL_TK[390] 
+ WL_TK[391] WL_TK[392] WL_TK[393] WL_TK[394] WL_TK[395] WL_TK[396] WL_TK[397] 
+ WL_TK[398] WL_TK[399] WL_TK[400] WL_TK[401] WL_TK[402] WL_TK[403] WL_TK[404] 
+ WL_TK[405] WL_TK[406] WL_TK[407] WL_TK[408] WL_TK[409] WL_TK[410] WL_TK[411] 
+ WL_TK[412] WL_TK[413] WL_TK[414] WL_TK[415] WL_TK[416] WL_TK[417] WL_TK[418] 
+ WL_TK[419] WL_TK[420] WL_TK[421] WL_TK[422] WL_TK[423] WL_TK[424] WL_TK[425] 
+ WL_TK[426] WL_TK[427] WL_TK[428] WL_TK[429] WL_TK[430] WL_TK[431] WL_TK[432] 
+ WL_TK[433] WL_TK[434] WL_TK[435] WL_TK[436] WL_TK[437] WL_TK[438] WL_TK[439] 
+ WL_TK[440] WL_TK[441] WL_TK[442] WL_TK[443] WL_TK[444] WL_TK[445] WL_TK[446] 
+ WL_TK[447] WL_TK[448] WL_TK[449] WL_TK[450] WL_TK[451] WL_TK[452] WL_TK[453] 
+ WL_TK[454] WL_TK[455] WL_TK[456] WL_TK[457] WL_TK[458] WL_TK[459] WL_TK[460] 
+ WL_TK[461] WL_TK[462] WL_TK[463] WL_TK[464] WL_TK[465] WL_TK[466] WL_TK[467] 
+ WL_TK[468] WL_TK[469] WL_TK[470] WL_TK[471] WL_TK[472] WL_TK[473] WL_TK[474] 
+ WL_TK[475] WL_TK[476] WL_TK[477] WL_TK[478] WL_TK[479] WL_TK[480] WL_TK[481] 
+ WL_TK[482] WL_TK[483] WL_TK[484] WL_TK[485] WL_TK[486] WL_TK[487] WL_TK[488] 
+ WL_TK[489] WL_TK[490] WL_TK[491] WL_TK[492] WL_TK[493] WL_TK[494] WL_TK[495] 
+ WL_TK[496] WL_TK[497] WL_TK[498] WL_TK[499] WL_TK[500] WL_TK[501] WL_TK[502] 
+ WL_TK[503] WL_TK[504] WL_TK[505] WL_TK[506] WL_TK[507] WL_TK[508] WL_TK[509] 
+ WL_TK[510] WL_TK[511] TIEH TIEL
*.PININFO BL_TK:B VDDI:B VSSI:B WL[0]:B WL[1]:B WL[2]:B WL[3]:B WL[4]:B 
*.PININFO WL[5]:B WL[6]:B WL[7]:B WL[8]:B WL[9]:B WL[10]:B WL[11]:B WL[12]:B 
*.PININFO WL[13]:B WL[14]:B WL[15]:B WL[16]:B WL[17]:B WL[18]:B WL[19]:B 
*.PININFO WL[20]:B WL[21]:B WL[22]:B WL[23]:B WL[24]:B WL[25]:B WL[26]:B 
*.PININFO WL[27]:B WL[28]:B WL[29]:B WL[30]:B WL[31]:B WL[32]:B WL[33]:B 
*.PININFO WL[34]:B WL[35]:B WL[36]:B WL[37]:B WL[38]:B WL[39]:B WL[40]:B 
*.PININFO WL[41]:B WL[42]:B WL[43]:B WL[44]:B WL[45]:B WL[46]:B WL[47]:B 
*.PININFO WL[48]:B WL[49]:B WL[50]:B WL[51]:B WL[52]:B WL[53]:B WL[54]:B 
*.PININFO WL[55]:B WL[56]:B WL[57]:B WL[58]:B WL[59]:B WL[60]:B WL[61]:B 
*.PININFO WL[62]:B WL[63]:B WL[64]:B WL[65]:B WL[66]:B WL[67]:B WL[68]:B 
*.PININFO WL[69]:B WL[70]:B WL[71]:B WL[72]:B WL[73]:B WL[74]:B WL[75]:B 
*.PININFO WL[76]:B WL[77]:B WL[78]:B WL[79]:B WL[80]:B WL[81]:B WL[82]:B 
*.PININFO WL[83]:B WL[84]:B WL[85]:B WL[86]:B WL[87]:B WL[88]:B WL[89]:B 
*.PININFO WL[90]:B WL[91]:B WL[92]:B WL[93]:B WL[94]:B WL[95]:B WL[96]:B 
*.PININFO WL[97]:B WL[98]:B WL[99]:B WL[100]:B WL[101]:B WL[102]:B WL[103]:B 
*.PININFO WL[104]:B WL[105]:B WL[106]:B WL[107]:B WL[108]:B WL[109]:B 
*.PININFO WL[110]:B WL[111]:B WL[112]:B WL[113]:B WL[114]:B WL[115]:B 
*.PININFO WL[116]:B WL[117]:B WL[118]:B WL[119]:B WL[120]:B WL[121]:B 
*.PININFO WL[122]:B WL[123]:B WL[124]:B WL[125]:B WL[126]:B WL[127]:B 
*.PININFO WL[128]:B WL[129]:B WL[130]:B WL[131]:B WL[132]:B WL[133]:B 
*.PININFO WL[134]:B WL[135]:B WL[136]:B WL[137]:B WL[138]:B WL[139]:B 
*.PININFO WL[140]:B WL[141]:B WL[142]:B WL[143]:B WL[144]:B WL[145]:B 
*.PININFO WL[146]:B WL[147]:B WL[148]:B WL[149]:B WL[150]:B WL[151]:B 
*.PININFO WL[152]:B WL[153]:B WL[154]:B WL[155]:B WL[156]:B WL[157]:B 
*.PININFO WL[158]:B WL[159]:B WL[160]:B WL[161]:B WL[162]:B WL[163]:B 
*.PININFO WL[164]:B WL[165]:B WL[166]:B WL[167]:B WL[168]:B WL[169]:B 
*.PININFO WL[170]:B WL[171]:B WL[172]:B WL[173]:B WL[174]:B WL[175]:B 
*.PININFO WL[176]:B WL[177]:B WL[178]:B WL[179]:B WL[180]:B WL[181]:B 
*.PININFO WL[182]:B WL[183]:B WL[184]:B WL[185]:B WL[186]:B WL[187]:B 
*.PININFO WL[188]:B WL[189]:B WL[190]:B WL[191]:B WL[192]:B WL[193]:B 
*.PININFO WL[194]:B WL[195]:B WL[196]:B WL[197]:B WL[198]:B WL[199]:B 
*.PININFO WL[200]:B WL[201]:B WL[202]:B WL[203]:B WL[204]:B WL[205]:B 
*.PININFO WL[206]:B WL[207]:B WL[208]:B WL[209]:B WL[210]:B WL[211]:B 
*.PININFO WL[212]:B WL[213]:B WL[214]:B WL[215]:B WL[216]:B WL[217]:B 
*.PININFO WL[218]:B WL[219]:B WL[220]:B WL[221]:B WL[222]:B WL[223]:B 
*.PININFO WL[224]:B WL[225]:B WL[226]:B WL[227]:B WL[228]:B WL[229]:B 
*.PININFO WL[230]:B WL[231]:B WL[232]:B WL[233]:B WL[234]:B WL[235]:B 
*.PININFO WL[236]:B WL[237]:B WL[238]:B WL[239]:B WL[240]:B WL[241]:B 
*.PININFO WL[242]:B WL[243]:B WL[244]:B WL[245]:B WL[246]:B WL[247]:B 
*.PININFO WL[248]:B WL[249]:B WL[250]:B WL[251]:B WL[252]:B WL[253]:B 
*.PININFO WL[254]:B WL[255]:B WL[256]:B WL[257]:B WL[258]:B WL[259]:B 
*.PININFO WL[260]:B WL[261]:B WL[262]:B WL[263]:B WL[264]:B WL[265]:B 
*.PININFO WL[266]:B WL[267]:B WL[268]:B WL[269]:B WL[270]:B WL[271]:B 
*.PININFO WL[272]:B WL[273]:B WL[274]:B WL[275]:B WL[276]:B WL[277]:B 
*.PININFO WL[278]:B WL[279]:B WL[280]:B WL[281]:B WL[282]:B WL[283]:B 
*.PININFO WL[284]:B WL[285]:B WL[286]:B WL[287]:B WL[288]:B WL[289]:B 
*.PININFO WL[290]:B WL[291]:B WL[292]:B WL[293]:B WL[294]:B WL[295]:B 
*.PININFO WL[296]:B WL[297]:B WL[298]:B WL[299]:B WL[300]:B WL[301]:B 
*.PININFO WL[302]:B WL[303]:B WL[304]:B WL[305]:B WL[306]:B WL[307]:B 
*.PININFO WL[308]:B WL[309]:B WL[310]:B WL[311]:B WL[312]:B WL[313]:B 
*.PININFO WL[314]:B WL[315]:B WL[316]:B WL[317]:B WL[318]:B WL[319]:B 
*.PININFO WL[320]:B WL[321]:B WL[322]:B WL[323]:B WL[324]:B WL[325]:B 
*.PININFO WL[326]:B WL[327]:B WL[328]:B WL[329]:B WL[330]:B WL[331]:B 
*.PININFO WL[332]:B WL[333]:B WL[334]:B WL[335]:B WL[336]:B WL[337]:B 
*.PININFO WL[338]:B WL[339]:B WL[340]:B WL[341]:B WL[342]:B WL[343]:B 
*.PININFO WL[344]:B WL[345]:B WL[346]:B WL[347]:B WL[348]:B WL[349]:B 
*.PININFO WL[350]:B WL[351]:B WL[352]:B WL[353]:B WL[354]:B WL[355]:B 
*.PININFO WL[356]:B WL[357]:B WL[358]:B WL[359]:B WL[360]:B WL[361]:B 
*.PININFO WL[362]:B WL[363]:B WL[364]:B WL[365]:B WL[366]:B WL[367]:B 
*.PININFO WL[368]:B WL[369]:B WL[370]:B WL[371]:B WL[372]:B WL[373]:B 
*.PININFO WL[374]:B WL[375]:B WL[376]:B WL[377]:B WL[378]:B WL[379]:B 
*.PININFO WL[380]:B WL[381]:B WL[382]:B WL[383]:B WL[384]:B WL[385]:B 
*.PININFO WL[386]:B WL[387]:B WL[388]:B WL[389]:B WL[390]:B WL[391]:B 
*.PININFO WL[392]:B WL[393]:B WL[394]:B WL[395]:B WL[396]:B WL[397]:B 
*.PININFO WL[398]:B WL[399]:B WL[400]:B WL[401]:B WL[402]:B WL[403]:B 
*.PININFO WL[404]:B WL[405]:B WL[406]:B WL[407]:B WL[408]:B WL[409]:B 
*.PININFO WL[410]:B WL[411]:B WL[412]:B WL[413]:B WL[414]:B WL[415]:B 
*.PININFO WL[416]:B WL[417]:B WL[418]:B WL[419]:B WL[420]:B WL[421]:B 
*.PININFO WL[422]:B WL[423]:B WL[424]:B WL[425]:B WL[426]:B WL[427]:B 
*.PININFO WL[428]:B WL[429]:B WL[430]:B WL[431]:B WL[432]:B WL[433]:B 
*.PININFO WL[434]:B WL[435]:B WL[436]:B WL[437]:B WL[438]:B WL[439]:B 
*.PININFO WL[440]:B WL[441]:B WL[442]:B WL[443]:B WL[444]:B WL[445]:B 
*.PININFO WL[446]:B WL[447]:B WL[448]:B WL[449]:B WL[450]:B WL[451]:B 
*.PININFO WL[452]:B WL[453]:B WL[454]:B WL[455]:B WL[456]:B WL[457]:B 
*.PININFO WL[458]:B WL[459]:B WL[460]:B WL[461]:B WL[462]:B WL[463]:B 
*.PININFO WL[464]:B WL[465]:B WL[466]:B WL[467]:B WL[468]:B WL[469]:B 
*.PININFO WL[470]:B WL[471]:B WL[472]:B WL[473]:B WL[474]:B WL[475]:B 
*.PININFO WL[476]:B WL[477]:B WL[478]:B WL[479]:B WL[480]:B WL[481]:B 
*.PININFO WL[482]:B WL[483]:B WL[484]:B WL[485]:B WL[486]:B WL[487]:B 
*.PININFO WL[488]:B WL[489]:B WL[490]:B WL[491]:B WL[492]:B WL[493]:B 
*.PININFO WL[494]:B WL[495]:B WL[496]:B WL[497]:B WL[498]:B WL[499]:B 
*.PININFO WL[500]:B WL[501]:B WL[502]:B WL[503]:B WL[504]:B WL[505]:B 
*.PININFO WL[506]:B WL[507]:B WL[508]:B WL[509]:B WL[510]:B WL[511]:B 
*.PININFO WL_TK[0]:B WL_TK[1]:B WL_TK[2]:B WL_TK[3]:B WL_TK[4]:B WL_TK[5]:B 
*.PININFO WL_TK[6]:B WL_TK[7]:B WL_TK[8]:B WL_TK[9]:B WL_TK[10]:B WL_TK[11]:B 
*.PININFO WL_TK[12]:B WL_TK[13]:B WL_TK[14]:B WL_TK[15]:B WL_TK[16]:B 
*.PININFO WL_TK[17]:B WL_TK[18]:B WL_TK[19]:B WL_TK[20]:B WL_TK[21]:B 
*.PININFO WL_TK[22]:B WL_TK[23]:B WL_TK[24]:B WL_TK[25]:B WL_TK[26]:B 
*.PININFO WL_TK[27]:B WL_TK[28]:B WL_TK[29]:B WL_TK[30]:B WL_TK[31]:B 
*.PININFO WL_TK[32]:B WL_TK[33]:B WL_TK[34]:B WL_TK[35]:B WL_TK[36]:B 
*.PININFO WL_TK[37]:B WL_TK[38]:B WL_TK[39]:B WL_TK[40]:B WL_TK[41]:B 
*.PININFO WL_TK[42]:B WL_TK[43]:B WL_TK[44]:B WL_TK[45]:B WL_TK[46]:B 
*.PININFO WL_TK[47]:B WL_TK[48]:B WL_TK[49]:B WL_TK[50]:B WL_TK[51]:B 
*.PININFO WL_TK[52]:B WL_TK[53]:B WL_TK[54]:B WL_TK[55]:B WL_TK[56]:B 
*.PININFO WL_TK[57]:B WL_TK[58]:B WL_TK[59]:B WL_TK[60]:B WL_TK[61]:B 
*.PININFO WL_TK[62]:B WL_TK[63]:B WL_TK[64]:B WL_TK[65]:B WL_TK[66]:B 
*.PININFO WL_TK[67]:B WL_TK[68]:B WL_TK[69]:B WL_TK[70]:B WL_TK[71]:B 
*.PININFO WL_TK[72]:B WL_TK[73]:B WL_TK[74]:B WL_TK[75]:B WL_TK[76]:B 
*.PININFO WL_TK[77]:B WL_TK[78]:B WL_TK[79]:B WL_TK[80]:B WL_TK[81]:B 
*.PININFO WL_TK[82]:B WL_TK[83]:B WL_TK[84]:B WL_TK[85]:B WL_TK[86]:B 
*.PININFO WL_TK[87]:B WL_TK[88]:B WL_TK[89]:B WL_TK[90]:B WL_TK[91]:B 
*.PININFO WL_TK[92]:B WL_TK[93]:B WL_TK[94]:B WL_TK[95]:B WL_TK[96]:B 
*.PININFO WL_TK[97]:B WL_TK[98]:B WL_TK[99]:B WL_TK[100]:B WL_TK[101]:B 
*.PININFO WL_TK[102]:B WL_TK[103]:B WL_TK[104]:B WL_TK[105]:B WL_TK[106]:B 
*.PININFO WL_TK[107]:B WL_TK[108]:B WL_TK[109]:B WL_TK[110]:B WL_TK[111]:B 
*.PININFO WL_TK[112]:B WL_TK[113]:B WL_TK[114]:B WL_TK[115]:B WL_TK[116]:B 
*.PININFO WL_TK[117]:B WL_TK[118]:B WL_TK[119]:B WL_TK[120]:B WL_TK[121]:B 
*.PININFO WL_TK[122]:B WL_TK[123]:B WL_TK[124]:B WL_TK[125]:B WL_TK[126]:B 
*.PININFO WL_TK[127]:B WL_TK[128]:B WL_TK[129]:B WL_TK[130]:B WL_TK[131]:B 
*.PININFO WL_TK[132]:B WL_TK[133]:B WL_TK[134]:B WL_TK[135]:B WL_TK[136]:B 
*.PININFO WL_TK[137]:B WL_TK[138]:B WL_TK[139]:B WL_TK[140]:B WL_TK[141]:B 
*.PININFO WL_TK[142]:B WL_TK[143]:B WL_TK[144]:B WL_TK[145]:B WL_TK[146]:B 
*.PININFO WL_TK[147]:B WL_TK[148]:B WL_TK[149]:B WL_TK[150]:B WL_TK[151]:B 
*.PININFO WL_TK[152]:B WL_TK[153]:B WL_TK[154]:B WL_TK[155]:B WL_TK[156]:B 
*.PININFO WL_TK[157]:B WL_TK[158]:B WL_TK[159]:B WL_TK[160]:B WL_TK[161]:B 
*.PININFO WL_TK[162]:B WL_TK[163]:B WL_TK[164]:B WL_TK[165]:B WL_TK[166]:B 
*.PININFO WL_TK[167]:B WL_TK[168]:B WL_TK[169]:B WL_TK[170]:B WL_TK[171]:B 
*.PININFO WL_TK[172]:B WL_TK[173]:B WL_TK[174]:B WL_TK[175]:B WL_TK[176]:B 
*.PININFO WL_TK[177]:B WL_TK[178]:B WL_TK[179]:B WL_TK[180]:B WL_TK[181]:B 
*.PININFO WL_TK[182]:B WL_TK[183]:B WL_TK[184]:B WL_TK[185]:B WL_TK[186]:B 
*.PININFO WL_TK[187]:B WL_TK[188]:B WL_TK[189]:B WL_TK[190]:B WL_TK[191]:B 
*.PININFO WL_TK[192]:B WL_TK[193]:B WL_TK[194]:B WL_TK[195]:B WL_TK[196]:B 
*.PININFO WL_TK[197]:B WL_TK[198]:B WL_TK[199]:B WL_TK[200]:B WL_TK[201]:B 
*.PININFO WL_TK[202]:B WL_TK[203]:B WL_TK[204]:B WL_TK[205]:B WL_TK[206]:B 
*.PININFO WL_TK[207]:B WL_TK[208]:B WL_TK[209]:B WL_TK[210]:B WL_TK[211]:B 
*.PININFO WL_TK[212]:B WL_TK[213]:B WL_TK[214]:B WL_TK[215]:B WL_TK[216]:B 
*.PININFO WL_TK[217]:B WL_TK[218]:B WL_TK[219]:B WL_TK[220]:B WL_TK[221]:B 
*.PININFO WL_TK[222]:B WL_TK[223]:B WL_TK[224]:B WL_TK[225]:B WL_TK[226]:B 
*.PININFO WL_TK[227]:B WL_TK[228]:B WL_TK[229]:B WL_TK[230]:B WL_TK[231]:B 
*.PININFO WL_TK[232]:B WL_TK[233]:B WL_TK[234]:B WL_TK[235]:B WL_TK[236]:B 
*.PININFO WL_TK[237]:B WL_TK[238]:B WL_TK[239]:B WL_TK[240]:B WL_TK[241]:B 
*.PININFO WL_TK[242]:B WL_TK[243]:B WL_TK[244]:B WL_TK[245]:B WL_TK[246]:B 
*.PININFO WL_TK[247]:B WL_TK[248]:B WL_TK[249]:B WL_TK[250]:B WL_TK[251]:B 
*.PININFO WL_TK[252]:B WL_TK[253]:B WL_TK[254]:B WL_TK[255]:B WL_TK[256]:B 
*.PININFO WL_TK[257]:B WL_TK[258]:B WL_TK[259]:B WL_TK[260]:B WL_TK[261]:B 
*.PININFO WL_TK[262]:B WL_TK[263]:B WL_TK[264]:B WL_TK[265]:B WL_TK[266]:B 
*.PININFO WL_TK[267]:B WL_TK[268]:B WL_TK[269]:B WL_TK[270]:B WL_TK[271]:B 
*.PININFO WL_TK[272]:B WL_TK[273]:B WL_TK[274]:B WL_TK[275]:B WL_TK[276]:B 
*.PININFO WL_TK[277]:B WL_TK[278]:B WL_TK[279]:B WL_TK[280]:B WL_TK[281]:B 
*.PININFO WL_TK[282]:B WL_TK[283]:B WL_TK[284]:B WL_TK[285]:B WL_TK[286]:B 
*.PININFO WL_TK[287]:B WL_TK[288]:B WL_TK[289]:B WL_TK[290]:B WL_TK[291]:B 
*.PININFO WL_TK[292]:B WL_TK[293]:B WL_TK[294]:B WL_TK[295]:B WL_TK[296]:B 
*.PININFO WL_TK[297]:B WL_TK[298]:B WL_TK[299]:B WL_TK[300]:B WL_TK[301]:B 
*.PININFO WL_TK[302]:B WL_TK[303]:B WL_TK[304]:B WL_TK[305]:B WL_TK[306]:B 
*.PININFO WL_TK[307]:B WL_TK[308]:B WL_TK[309]:B WL_TK[310]:B WL_TK[311]:B 
*.PININFO WL_TK[312]:B WL_TK[313]:B WL_TK[314]:B WL_TK[315]:B WL_TK[316]:B 
*.PININFO WL_TK[317]:B WL_TK[318]:B WL_TK[319]:B WL_TK[320]:B WL_TK[321]:B 
*.PININFO WL_TK[322]:B WL_TK[323]:B WL_TK[324]:B WL_TK[325]:B WL_TK[326]:B 
*.PININFO WL_TK[327]:B WL_TK[328]:B WL_TK[329]:B WL_TK[330]:B WL_TK[331]:B 
*.PININFO WL_TK[332]:B WL_TK[333]:B WL_TK[334]:B WL_TK[335]:B WL_TK[336]:B 
*.PININFO WL_TK[337]:B WL_TK[338]:B WL_TK[339]:B WL_TK[340]:B WL_TK[341]:B 
*.PININFO WL_TK[342]:B WL_TK[343]:B WL_TK[344]:B WL_TK[345]:B WL_TK[346]:B 
*.PININFO WL_TK[347]:B WL_TK[348]:B WL_TK[349]:B WL_TK[350]:B WL_TK[351]:B 
*.PININFO WL_TK[352]:B WL_TK[353]:B WL_TK[354]:B WL_TK[355]:B WL_TK[356]:B 
*.PININFO WL_TK[357]:B WL_TK[358]:B WL_TK[359]:B WL_TK[360]:B WL_TK[361]:B 
*.PININFO WL_TK[362]:B WL_TK[363]:B WL_TK[364]:B WL_TK[365]:B WL_TK[366]:B 
*.PININFO WL_TK[367]:B WL_TK[368]:B WL_TK[369]:B WL_TK[370]:B WL_TK[371]:B 
*.PININFO WL_TK[372]:B WL_TK[373]:B WL_TK[374]:B WL_TK[375]:B WL_TK[376]:B 
*.PININFO WL_TK[377]:B WL_TK[378]:B WL_TK[379]:B WL_TK[380]:B WL_TK[381]:B 
*.PININFO WL_TK[382]:B WL_TK[383]:B WL_TK[384]:B WL_TK[385]:B WL_TK[386]:B 
*.PININFO WL_TK[387]:B WL_TK[388]:B WL_TK[389]:B WL_TK[390]:B WL_TK[391]:B 
*.PININFO WL_TK[392]:B WL_TK[393]:B WL_TK[394]:B WL_TK[395]:B WL_TK[396]:B 
*.PININFO WL_TK[397]:B WL_TK[398]:B WL_TK[399]:B WL_TK[400]:B WL_TK[401]:B 
*.PININFO WL_TK[402]:B WL_TK[403]:B WL_TK[404]:B WL_TK[405]:B WL_TK[406]:B 
*.PININFO WL_TK[407]:B WL_TK[408]:B WL_TK[409]:B WL_TK[410]:B WL_TK[411]:B 
*.PININFO WL_TK[412]:B WL_TK[413]:B WL_TK[414]:B WL_TK[415]:B WL_TK[416]:B 
*.PININFO WL_TK[417]:B WL_TK[418]:B WL_TK[419]:B WL_TK[420]:B WL_TK[421]:B 
*.PININFO WL_TK[422]:B WL_TK[423]:B WL_TK[424]:B WL_TK[425]:B WL_TK[426]:B 
*.PININFO WL_TK[427]:B WL_TK[428]:B WL_TK[429]:B WL_TK[430]:B WL_TK[431]:B 
*.PININFO WL_TK[432]:B WL_TK[433]:B WL_TK[434]:B WL_TK[435]:B WL_TK[436]:B 
*.PININFO WL_TK[437]:B WL_TK[438]:B WL_TK[439]:B WL_TK[440]:B WL_TK[441]:B 
*.PININFO WL_TK[442]:B WL_TK[443]:B WL_TK[444]:B WL_TK[445]:B WL_TK[446]:B 
*.PININFO WL_TK[447]:B WL_TK[448]:B WL_TK[449]:B WL_TK[450]:B WL_TK[451]:B 
*.PININFO WL_TK[452]:B WL_TK[453]:B WL_TK[454]:B WL_TK[455]:B WL_TK[456]:B 
*.PININFO WL_TK[457]:B WL_TK[458]:B WL_TK[459]:B WL_TK[460]:B WL_TK[461]:B 
*.PININFO WL_TK[462]:B WL_TK[463]:B WL_TK[464]:B WL_TK[465]:B WL_TK[466]:B 
*.PININFO WL_TK[467]:B WL_TK[468]:B WL_TK[469]:B WL_TK[470]:B WL_TK[471]:B 
*.PININFO WL_TK[472]:B WL_TK[473]:B WL_TK[474]:B WL_TK[475]:B WL_TK[476]:B 
*.PININFO WL_TK[477]:B WL_TK[478]:B WL_TK[479]:B WL_TK[480]:B WL_TK[481]:B 
*.PININFO WL_TK[482]:B WL_TK[483]:B WL_TK[484]:B WL_TK[485]:B WL_TK[486]:B 
*.PININFO WL_TK[487]:B WL_TK[488]:B WL_TK[489]:B WL_TK[490]:B WL_TK[491]:B 
*.PININFO WL_TK[492]:B WL_TK[493]:B WL_TK[494]:B WL_TK[495]:B WL_TK[496]:B 
*.PININFO WL_TK[497]:B WL_TK[498]:B WL_TK[499]:B WL_TK[500]:B WL_TK[501]:B 
*.PININFO WL_TK[502]:B WL_TK[503]:B WL_TK[504]:B WL_TK[505]:B WL_TK[506]:B 
*.PININFO WL_TK[507]:B WL_TK[508]:B WL_TK[509]:B WL_TK[510]:B WL_TK[511]:B 
*.PININFO TIEH:B TIEL:B
XTRKNORX64_DUMY6 BL_TK VDDI VSSI WL[256] WL[257] WL[258] WL[259] WL[260] 
+ WL[261] WL[262] WL[263] WL[264] WL[265] WL[266] WL[267] WL[268] WL[269] 
+ WL[270] WL[271] WL[272] WL[273] WL[274] WL[275] WL[276] WL[277] WL[278] 
+ WL[279] WL[280] WL[281] WL[282] WL[283] WL[284] WL[285] WL[286] WL[287] 
+ WL[288] WL[289] WL[290] WL[291] WL[292] WL[293] WL[294] WL[295] WL[296] 
+ WL[297] WL[298] WL[299] WL[300] WL[301] WL[302] WL[303] WL[304] WL[305] 
+ WL[306] WL[307] WL[308] WL[309] WL[310] WL[311] WL[312] WL[313] WL[314] 
+ WL[315] WL[316] WL[317] WL[318] WL[319] WL_TK[256] WL_TK[257] WL_TK[258] 
+ WL_TK[259] WL_TK[260] WL_TK[261] WL_TK[262] WL_TK[263] WL_TK[264] WL_TK[265] 
+ WL_TK[266] WL_TK[267] WL_TK[268] WL_TK[269] WL_TK[270] WL_TK[271] WL_TK[272] 
+ WL_TK[273] WL_TK[274] WL_TK[275] WL_TK[276] WL_TK[277] WL_TK[278] WL_TK[279] 
+ WL_TK[280] WL_TK[281] WL_TK[282] WL_TK[283] WL_TK[284] WL_TK[285] WL_TK[286] 
+ WL_TK[287] WL_TK[288] WL_TK[289] WL_TK[290] WL_TK[291] WL_TK[292] WL_TK[293] 
+ WL_TK[294] WL_TK[295] WL_TK[296] WL_TK[297] WL_TK[298] WL_TK[299] WL_TK[300] 
+ WL_TK[301] WL_TK[302] WL_TK[303] WL_TK[304] WL_TK[305] WL_TK[306] WL_TK[307] 
+ WL_TK[308] WL_TK[309] WL_TK[310] WL_TK[311] WL_TK[312] WL_TK[313] WL_TK[314] 
+ WL_TK[315] WL_TK[316] WL_TK[317] WL_TK[318] WL_TK[319] NET49[0] NET49[1] 
+ NET49[2] NET49[3] NET49[4] NET49[5] NET49[6] NET49[7] NET49[8] NET49[9] 
+ NET49[10] NET49[11] NET49[12] NET49[13] NET49[14] NET49[15] NET49[16] 
+ NET49[17] NET49[18] NET49[19] NET49[20] NET49[21] NET49[22] NET49[23] 
+ NET49[24] NET49[25] NET49[26] NET49[27] NET49[28] NET49[29] NET49[30] 
+ NET49[31] NET48 NET47 NET46[0] NET46[1] NET46[2] NET46[3] NET46[4] NET46[5] 
+ NET46[6] NET46[7] NET46[8] NET46[9] NET46[10] NET46[11] NET46[12] NET46[13] 
+ NET46[14] NET46[15] NET46[16] NET46[17] NET46[18] NET46[19] NET46[20] 
+ NET46[21] NET46[22] NET46[23] NET46[24] NET46[25] NET46[26] NET46[27] 
+ NET46[28] NET46[29] NET46[30] NET46[31] TIEH S1AHSF400W40_TRKNORX64_CHAR
XTRKNORX64_DUMY4 BL_TK VDDI VSSI WL[128] WL[129] WL[130] WL[131] WL[132] 
+ WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] WL[140] WL[141] 
+ WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] WL[149] WL[150] 
+ WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] WL[158] WL[159] 
+ WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] WL[167] WL[168] 
+ WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] WL[176] WL[177] 
+ WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] WL[185] WL[186] 
+ WL[187] WL[188] WL[189] WL[190] WL[191] WL_TK[128] WL_TK[129] WL_TK[130] 
+ WL_TK[131] WL_TK[132] WL_TK[133] WL_TK[134] WL_TK[135] WL_TK[136] WL_TK[137] 
+ WL_TK[138] WL_TK[139] WL_TK[140] WL_TK[141] WL_TK[142] WL_TK[143] WL_TK[144] 
+ WL_TK[145] WL_TK[146] WL_TK[147] WL_TK[148] WL_TK[149] WL_TK[150] WL_TK[151] 
+ WL_TK[152] WL_TK[153] WL_TK[154] WL_TK[155] WL_TK[156] WL_TK[157] WL_TK[158] 
+ WL_TK[159] WL_TK[160] WL_TK[161] WL_TK[162] WL_TK[163] WL_TK[164] WL_TK[165] 
+ WL_TK[166] WL_TK[167] WL_TK[168] WL_TK[169] WL_TK[170] WL_TK[171] WL_TK[172] 
+ WL_TK[173] WL_TK[174] WL_TK[175] WL_TK[176] WL_TK[177] WL_TK[178] WL_TK[179] 
+ WL_TK[180] WL_TK[181] WL_TK[182] WL_TK[183] WL_TK[184] WL_TK[185] WL_TK[186] 
+ WL_TK[187] WL_TK[188] WL_TK[189] WL_TK[190] WL_TK[191] NET59[0] NET59[1] 
+ NET59[2] NET59[3] NET59[4] NET59[5] NET59[6] NET59[7] NET59[8] NET59[9] 
+ NET59[10] NET59[11] NET59[12] NET59[13] NET59[14] NET59[15] NET59[16] 
+ NET59[17] NET59[18] NET59[19] NET59[20] NET59[21] NET59[22] NET59[23] 
+ NET59[24] NET59[25] NET59[26] NET59[27] NET59[28] NET59[29] NET59[30] 
+ NET59[31] NET58 NET57 NET56[0] NET56[1] NET56[2] NET56[3] NET56[4] NET56[5] 
+ NET56[6] NET56[7] NET56[8] NET56[9] NET56[10] NET56[11] NET56[12] NET56[13] 
+ NET56[14] NET56[15] NET56[16] NET56[17] NET56[18] NET56[19] NET56[20] 
+ NET56[21] NET56[22] NET56[23] NET56[24] NET56[25] NET56[26] NET56[27] 
+ NET56[28] NET56[29] NET56[30] NET56[31] TIEH S1AHSF400W40_TRKNORX64_CHAR
XTRKNORX64_DUMY7 BL_TK VDDI VSSI WL[320] WL[321] WL[322] WL[323] WL[324] 
+ WL[325] WL[326] WL[327] WL[328] WL[329] WL[330] WL[331] WL[332] WL[333] 
+ WL[334] WL[335] WL[336] WL[337] WL[338] WL[339] WL[340] WL[341] WL[342] 
+ WL[343] WL[344] WL[345] WL[346] WL[347] WL[348] WL[349] WL[350] WL[351] 
+ WL[352] WL[353] WL[354] WL[355] WL[356] WL[357] WL[358] WL[359] WL[360] 
+ WL[361] WL[362] WL[363] WL[364] WL[365] WL[366] WL[367] WL[368] WL[369] 
+ WL[370] WL[371] WL[372] WL[373] WL[374] WL[375] WL[376] WL[377] WL[378] 
+ WL[379] WL[380] WL[381] WL[382] WL[383] WL_TK[320] WL_TK[321] WL_TK[322] 
+ WL_TK[323] WL_TK[324] WL_TK[325] WL_TK[326] WL_TK[327] WL_TK[328] WL_TK[329] 
+ WL_TK[330] WL_TK[331] WL_TK[332] WL_TK[333] WL_TK[334] WL_TK[335] WL_TK[336] 
+ WL_TK[337] WL_TK[338] WL_TK[339] WL_TK[340] WL_TK[341] WL_TK[342] WL_TK[343] 
+ WL_TK[344] WL_TK[345] WL_TK[346] WL_TK[347] WL_TK[348] WL_TK[349] WL_TK[350] 
+ WL_TK[351] WL_TK[352] WL_TK[353] WL_TK[354] WL_TK[355] WL_TK[356] WL_TK[357] 
+ WL_TK[358] WL_TK[359] WL_TK[360] WL_TK[361] WL_TK[362] WL_TK[363] WL_TK[364] 
+ WL_TK[365] WL_TK[366] WL_TK[367] WL_TK[368] WL_TK[369] WL_TK[370] WL_TK[371] 
+ WL_TK[372] WL_TK[373] WL_TK[374] WL_TK[375] WL_TK[376] WL_TK[377] WL_TK[378] 
+ WL_TK[379] WL_TK[380] WL_TK[381] WL_TK[382] WL_TK[383] NET39[0] NET39[1] 
+ NET39[2] NET39[3] NET39[4] NET39[5] NET39[6] NET39[7] NET39[8] NET39[9] 
+ NET39[10] NET39[11] NET39[12] NET39[13] NET39[14] NET39[15] NET39[16] 
+ NET39[17] NET39[18] NET39[19] NET39[20] NET39[21] NET39[22] NET39[23] 
+ NET39[24] NET39[25] NET39[26] NET39[27] NET39[28] NET39[29] NET39[30] 
+ NET39[31] NET38 NET37 NET36[0] NET36[1] NET36[2] NET36[3] NET36[4] NET36[5] 
+ NET36[6] NET36[7] NET36[8] NET36[9] NET36[10] NET36[11] NET36[12] NET36[13] 
+ NET36[14] NET36[15] NET36[16] NET36[17] NET36[18] NET36[19] NET36[20] 
+ NET36[21] NET36[22] NET36[23] NET36[24] NET36[25] NET36[26] NET36[27] 
+ NET36[28] NET36[29] NET36[30] NET36[31] TIEH S1AHSF400W40_TRKNORX64_CHAR
XTRKNORX64_DUMY8 BL_TK VDDI VSSI WL[384] WL[385] WL[386] WL[387] WL[388] 
+ WL[389] WL[390] WL[391] WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] 
+ WL[398] WL[399] WL[400] WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] 
+ WL[407] WL[408] WL[409] WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] 
+ WL[416] WL[417] WL[418] WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] 
+ WL[425] WL[426] WL[427] WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] 
+ WL[434] WL[435] WL[436] WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] 
+ WL[443] WL[444] WL[445] WL[446] WL[447] WL_TK[384] WL_TK[385] WL_TK[386] 
+ WL_TK[387] WL_TK[388] WL_TK[389] WL_TK[390] WL_TK[391] WL_TK[392] WL_TK[393] 
+ WL_TK[394] WL_TK[395] WL_TK[396] WL_TK[397] WL_TK[398] WL_TK[399] WL_TK[400] 
+ WL_TK[401] WL_TK[402] WL_TK[403] WL_TK[404] WL_TK[405] WL_TK[406] WL_TK[407] 
+ WL_TK[408] WL_TK[409] WL_TK[410] WL_TK[411] WL_TK[412] WL_TK[413] WL_TK[414] 
+ WL_TK[415] WL_TK[416] WL_TK[417] WL_TK[418] WL_TK[419] WL_TK[420] WL_TK[421] 
+ WL_TK[422] WL_TK[423] WL_TK[424] WL_TK[425] WL_TK[426] WL_TK[427] WL_TK[428] 
+ WL_TK[429] WL_TK[430] WL_TK[431] WL_TK[432] WL_TK[433] WL_TK[434] WL_TK[435] 
+ WL_TK[436] WL_TK[437] WL_TK[438] WL_TK[439] WL_TK[440] WL_TK[441] WL_TK[442] 
+ WL_TK[443] WL_TK[444] WL_TK[445] WL_TK[446] WL_TK[447] NET29[0] NET29[1] 
+ NET29[2] NET29[3] NET29[4] NET29[5] NET29[6] NET29[7] NET29[8] NET29[9] 
+ NET29[10] NET29[11] NET29[12] NET29[13] NET29[14] NET29[15] NET29[16] 
+ NET29[17] NET29[18] NET29[19] NET29[20] NET29[21] NET29[22] NET29[23] 
+ NET29[24] NET29[25] NET29[26] NET29[27] NET29[28] NET29[29] NET29[30] 
+ NET29[31] NET28 NET27 NET26[0] NET26[1] NET26[2] NET26[3] NET26[4] NET26[5] 
+ NET26[6] NET26[7] NET26[8] NET26[9] NET26[10] NET26[11] NET26[12] NET26[13] 
+ NET26[14] NET26[15] NET26[16] NET26[17] NET26[18] NET26[19] NET26[20] 
+ NET26[21] NET26[22] NET26[23] NET26[24] NET26[25] NET26[26] NET26[27] 
+ NET26[28] NET26[29] NET26[30] NET26[31] TIEH S1AHSF400W40_TRKNORX64_CHAR
XTRKNORX64_DUMY9 BL_TK VDDI VSSI WL[448] WL[449] WL[450] WL[451] WL[452] 
+ WL[453] WL[454] WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] 
+ WL[462] WL[463] WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] 
+ WL[471] WL[472] WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] 
+ WL[480] WL[481] WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] 
+ WL[489] WL[490] WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] 
+ WL[498] WL[499] WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] 
+ WL[507] WL[508] WL[509] WL[510] WL[511] WL_TK[448] WL_TK[449] WL_TK[450] 
+ WL_TK[451] WL_TK[452] WL_TK[453] WL_TK[454] WL_TK[455] WL_TK[456] WL_TK[457] 
+ WL_TK[458] WL_TK[459] WL_TK[460] WL_TK[461] WL_TK[462] WL_TK[463] WL_TK[464] 
+ WL_TK[465] WL_TK[466] WL_TK[467] WL_TK[468] WL_TK[469] WL_TK[470] WL_TK[471] 
+ WL_TK[472] WL_TK[473] WL_TK[474] WL_TK[475] WL_TK[476] WL_TK[477] WL_TK[478] 
+ WL_TK[479] WL_TK[480] WL_TK[481] WL_TK[482] WL_TK[483] WL_TK[484] WL_TK[485] 
+ WL_TK[486] WL_TK[487] WL_TK[488] WL_TK[489] WL_TK[490] WL_TK[491] WL_TK[492] 
+ WL_TK[493] WL_TK[494] WL_TK[495] WL_TK[496] WL_TK[497] WL_TK[498] WL_TK[499] 
+ WL_TK[500] WL_TK[501] WL_TK[502] WL_TK[503] WL_TK[504] WL_TK[505] WL_TK[506] 
+ WL_TK[507] WL_TK[508] WL_TK[509] WL_TK[510] WL_TK[511] NET19[0] NET19[1] 
+ NET19[2] NET19[3] NET19[4] NET19[5] NET19[6] NET19[7] NET19[8] NET19[9] 
+ NET19[10] NET19[11] NET19[12] NET19[13] NET19[14] NET19[15] NET19[16] 
+ NET19[17] NET19[18] NET19[19] NET19[20] NET19[21] NET19[22] NET19[23] 
+ NET19[24] NET19[25] NET19[26] NET19[27] NET19[28] NET19[29] NET19[30] 
+ NET19[31] NET18 NET17 NET16[0] NET16[1] NET16[2] NET16[3] NET16[4] NET16[5] 
+ NET16[6] NET16[7] NET16[8] NET16[9] NET16[10] NET16[11] NET16[12] NET16[13] 
+ NET16[14] NET16[15] NET16[16] NET16[17] NET16[18] NET16[19] NET16[20] 
+ NET16[21] NET16[22] NET16[23] NET16[24] NET16[25] NET16[26] NET16[27] 
+ NET16[28] NET16[29] NET16[30] NET16[31] TIEH S1AHSF400W40_TRKNORX64_CHAR
XTRKNORX64_DUMY3 BL_TK VDDI VSSI WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] 
+ WL[70] WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] 
+ WL[81] WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] 
+ WL[92] WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] 
+ WL[102] WL[103] WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] 
+ WL[111] WL[112] WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] 
+ WL[120] WL[121] WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL_TK[64] 
+ WL_TK[65] WL_TK[66] WL_TK[67] WL_TK[68] WL_TK[69] WL_TK[70] WL_TK[71] 
+ WL_TK[72] WL_TK[73] WL_TK[74] WL_TK[75] WL_TK[76] WL_TK[77] WL_TK[78] 
+ WL_TK[79] WL_TK[80] WL_TK[81] WL_TK[82] WL_TK[83] WL_TK[84] WL_TK[85] 
+ WL_TK[86] WL_TK[87] WL_TK[88] WL_TK[89] WL_TK[90] WL_TK[91] WL_TK[92] 
+ WL_TK[93] WL_TK[94] WL_TK[95] WL_TK[96] WL_TK[97] WL_TK[98] WL_TK[99] 
+ WL_TK[100] WL_TK[101] WL_TK[102] WL_TK[103] WL_TK[104] WL_TK[105] WL_TK[106] 
+ WL_TK[107] WL_TK[108] WL_TK[109] WL_TK[110] WL_TK[111] WL_TK[112] WL_TK[113] 
+ WL_TK[114] WL_TK[115] WL_TK[116] WL_TK[117] WL_TK[118] WL_TK[119] WL_TK[120] 
+ WL_TK[121] WL_TK[122] WL_TK[123] WL_TK[124] WL_TK[125] WL_TK[126] WL_TK[127] 
+ NET69[0] NET69[1] NET69[2] NET69[3] NET69[4] NET69[5] NET69[6] NET69[7] 
+ NET69[8] NET69[9] NET69[10] NET69[11] NET69[12] NET69[13] NET69[14] 
+ NET69[15] NET69[16] NET69[17] NET69[18] NET69[19] NET69[20] NET69[21] 
+ NET69[22] NET69[23] NET69[24] NET69[25] NET69[26] NET69[27] NET69[28] 
+ NET69[29] NET69[30] NET69[31] NET68 NET67 NET66[0] NET66[1] NET66[2] 
+ NET66[3] NET66[4] NET66[5] NET66[6] NET66[7] NET66[8] NET66[9] NET66[10] 
+ NET66[11] NET66[12] NET66[13] NET66[14] NET66[15] NET66[16] NET66[17] 
+ NET66[18] NET66[19] NET66[20] NET66[21] NET66[22] NET66[23] NET66[24] 
+ NET66[25] NET66[26] NET66[27] NET66[28] NET66[29] NET66[30] NET66[31] TIEH 
+ S1AHSF400W40_TRKNORX64_CHAR
XTRKNORX64_DYMY5 BL_TK VDDI VSSI WL[192] WL[193] WL[194] WL[195] WL[196] 
+ WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] WL[203] WL[204] WL[205] 
+ WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] WL[212] WL[213] WL[214] 
+ WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] WL[221] WL[222] WL[223] 
+ WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] WL[230] WL[231] WL[232] 
+ WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] WL[239] WL[240] WL[241] 
+ WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] WL[248] WL[249] WL[250] 
+ WL[251] WL[252] WL[253] WL[254] WL[255] WL_TK[192] WL_TK[193] WL_TK[194] 
+ WL_TK[195] WL_TK[196] WL_TK[197] WL_TK[198] WL_TK[199] WL_TK[200] WL_TK[201] 
+ WL_TK[202] WL_TK[203] WL_TK[204] WL_TK[205] WL_TK[206] WL_TK[207] WL_TK[208] 
+ WL_TK[209] WL_TK[210] WL_TK[211] WL_TK[212] WL_TK[213] WL_TK[214] WL_TK[215] 
+ WL_TK[216] WL_TK[217] WL_TK[218] WL_TK[219] WL_TK[220] WL_TK[221] WL_TK[222] 
+ WL_TK[223] WL_TK[224] WL_TK[225] WL_TK[226] WL_TK[227] WL_TK[228] WL_TK[229] 
+ WL_TK[230] WL_TK[231] WL_TK[232] WL_TK[233] WL_TK[234] WL_TK[235] WL_TK[236] 
+ WL_TK[237] WL_TK[238] WL_TK[239] WL_TK[240] WL_TK[241] WL_TK[242] WL_TK[243] 
+ WL_TK[244] WL_TK[245] WL_TK[246] WL_TK[247] WL_TK[248] WL_TK[249] WL_TK[250] 
+ WL_TK[251] WL_TK[252] WL_TK[253] WL_TK[254] WL_TK[255] NET79[0] NET79[1] 
+ NET79[2] NET79[3] NET79[4] NET79[5] NET79[6] NET79[7] NET79[8] NET79[9] 
+ NET79[10] NET79[11] NET79[12] NET79[13] NET79[14] NET79[15] NET79[16] 
+ NET79[17] NET79[18] NET79[19] NET79[20] NET79[21] NET79[22] NET79[23] 
+ NET79[24] NET79[25] NET79[26] NET79[27] NET79[28] NET79[29] NET79[30] 
+ NET79[31] NET78 NET77 NET76[0] NET76[1] NET76[2] NET76[3] NET76[4] NET76[5] 
+ NET76[6] NET76[7] NET76[8] NET76[9] NET76[10] NET76[11] NET76[12] NET76[13] 
+ NET76[14] NET76[15] NET76[16] NET76[17] NET76[18] NET76[19] NET76[20] 
+ NET76[21] NET76[22] NET76[23] NET76[24] NET76[25] NET76[26] NET76[27] 
+ NET76[28] NET76[29] NET76[30] NET76[31] TIEH S1AHSF400W40_TRKNORX64_CHAR
XTRKNORX16_DUMY0 BL_TK VDDI VSSI WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] 
+ WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] 
+ WL_TK[16] WL_TK[17] WL_TK[18] WL_TK[19] WL_TK[20] WL_TK[21] WL_TK[22] 
+ WL_TK[23] WL_TK[24] WL_TK[25] WL_TK[26] WL_TK[27] WL_TK[28] WL_TK[29] 
+ WL_TK[30] WL_TK[31] NET89[0] NET89[1] NET89[2] NET89[3] NET89[4] NET89[5] 
+ NET89[6] NET89[7] NET88 NET108 NET86[0] NET86[1] NET86[2] NET86[3] NET86[4] 
+ NET86[5] NET86[6] NET86[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
XTRKNORX16_DUMY1 BL_TK VDDI VSSI WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] 
+ WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] 
+ WL_TK[32] WL_TK[33] WL_TK[34] WL_TK[35] WL_TK[36] WL_TK[37] WL_TK[38] 
+ WL_TK[39] WL_TK[40] WL_TK[41] WL_TK[42] WL_TK[43] WL_TK[44] WL_TK[45] 
+ WL_TK[46] WL_TK[47] NET99[0] NET99[1] NET99[2] NET99[3] NET99[4] NET99[5] 
+ NET99[6] NET99[7] NET98 NET88 NET96[0] NET96[1] NET96[2] NET96[3] NET96[4] 
+ NET96[5] NET96[6] NET96[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
XTRKNORX16_BCELL BL_TK VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] 
+ WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL_TK[0] 
+ WL_TK[1] WL_TK[2] WL_TK[3] WL_TK[4] WL_TK[5] WL_TK[6] WL_TK[7] WL_TK[8] 
+ WL_TK[9] WL_TK[10] WL_TK[11] WL_TK[12] WL_TK[13] WL_TK[14] WL_TK[15] 
+ NET109[0] NET109[1] NET109[2] NET109[3] NET109[4] NET109[5] NET109[6] 
+ NET109[7] NET108 NET107 NET106[0] NET106[1] NET106[2] NET106[3] NET106[4] 
+ NET106[5] NET106[6] NET106[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
XTRKNORX16_DUMY2 BL_TK VDDI VSSI WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] 
+ WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] 
+ WL_TK[48] WL_TK[49] WL_TK[50] WL_TK[51] WL_TK[52] WL_TK[53] WL_TK[54] 
+ WL_TK[55] WL_TK[56] WL_TK[57] WL_TK[58] WL_TK[59] WL_TK[60] WL_TK[61] 
+ WL_TK[62] WL_TK[63] NET119[0] NET119[1] NET119[2] NET119[3] NET119[4] 
+ NET119[5] NET119[6] NET119[7] NET118 NET98 NET116[0] NET116[1] NET116[2] 
+ NET116[3] NET116[4] NET116[5] NET116[6] NET116[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    TKBL_S64_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TKBL_S64_CHAR BL_TK VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL_TK[0] WL_TK[1] WL_TK[2] WL_TK[3] WL_TK[4] WL_TK[5] 
+ WL_TK[6] WL_TK[7] WL_TK[8] WL_TK[9] WL_TK[10] WL_TK[11] WL_TK[12] WL_TK[13] 
+ WL_TK[14] WL_TK[15] WL_TK[16] WL_TK[17] WL_TK[18] WL_TK[19] WL_TK[20] 
+ WL_TK[21] WL_TK[22] WL_TK[23] WL_TK[24] WL_TK[25] WL_TK[26] WL_TK[27] 
+ WL_TK[28] WL_TK[29] WL_TK[30] WL_TK[31] WL_TK[32] WL_TK[33] WL_TK[34] 
+ WL_TK[35] WL_TK[36] WL_TK[37] WL_TK[38] WL_TK[39] WL_TK[40] WL_TK[41] 
+ WL_TK[42] WL_TK[43] WL_TK[44] WL_TK[45] WL_TK[46] WL_TK[47] WL_TK[48] 
+ WL_TK[49] WL_TK[50] WL_TK[51] WL_TK[52] WL_TK[53] WL_TK[54] WL_TK[55] 
+ WL_TK[56] WL_TK[57] WL_TK[58] WL_TK[59] WL_TK[60] WL_TK[61] WL_TK[62] 
+ WL_TK[63] TIEH TIEL
*.PININFO BL_TK:B VDDI:B VSSI:B WL[0]:B WL[1]:B WL[2]:B WL[3]:B WL[4]:B 
*.PININFO WL[5]:B WL[6]:B WL[7]:B WL[8]:B WL[9]:B WL[10]:B WL[11]:B WL[12]:B 
*.PININFO WL[13]:B WL[14]:B WL[15]:B WL[16]:B WL[17]:B WL[18]:B WL[19]:B 
*.PININFO WL[20]:B WL[21]:B WL[22]:B WL[23]:B WL[24]:B WL[25]:B WL[26]:B 
*.PININFO WL[27]:B WL[28]:B WL[29]:B WL[30]:B WL[31]:B WL[32]:B WL[33]:B 
*.PININFO WL[34]:B WL[35]:B WL[36]:B WL[37]:B WL[38]:B WL[39]:B WL[40]:B 
*.PININFO WL[41]:B WL[42]:B WL[43]:B WL[44]:B WL[45]:B WL[46]:B WL[47]:B 
*.PININFO WL[48]:B WL[49]:B WL[50]:B WL[51]:B WL[52]:B WL[53]:B WL[54]:B 
*.PININFO WL[55]:B WL[56]:B WL[57]:B WL[58]:B WL[59]:B WL[60]:B WL[61]:B 
*.PININFO WL[62]:B WL[63]:B WL_TK[0]:B WL_TK[1]:B WL_TK[2]:B WL_TK[3]:B 
*.PININFO WL_TK[4]:B WL_TK[5]:B WL_TK[6]:B WL_TK[7]:B WL_TK[8]:B WL_TK[9]:B 
*.PININFO WL_TK[10]:B WL_TK[11]:B WL_TK[12]:B WL_TK[13]:B WL_TK[14]:B 
*.PININFO WL_TK[15]:B WL_TK[16]:B WL_TK[17]:B WL_TK[18]:B WL_TK[19]:B 
*.PININFO WL_TK[20]:B WL_TK[21]:B WL_TK[22]:B WL_TK[23]:B WL_TK[24]:B 
*.PININFO WL_TK[25]:B WL_TK[26]:B WL_TK[27]:B WL_TK[28]:B WL_TK[29]:B 
*.PININFO WL_TK[30]:B WL_TK[31]:B WL_TK[32]:B WL_TK[33]:B WL_TK[34]:B 
*.PININFO WL_TK[35]:B WL_TK[36]:B WL_TK[37]:B WL_TK[38]:B WL_TK[39]:B 
*.PININFO WL_TK[40]:B WL_TK[41]:B WL_TK[42]:B WL_TK[43]:B WL_TK[44]:B 
*.PININFO WL_TK[45]:B WL_TK[46]:B WL_TK[47]:B WL_TK[48]:B WL_TK[49]:B 
*.PININFO WL_TK[50]:B WL_TK[51]:B WL_TK[52]:B WL_TK[53]:B WL_TK[54]:B 
*.PININFO WL_TK[55]:B WL_TK[56]:B WL_TK[57]:B WL_TK[58]:B WL_TK[59]:B 
*.PININFO WL_TK[60]:B WL_TK[61]:B WL_TK[62]:B WL_TK[63]:B TIEH:B TIEL:B
XTRKNORX16_DUMY0 BL_TK VDDI VSSI WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] 
+ WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] 
+ WL_TK[16] WL_TK[17] WL_TK[18] WL_TK[19] WL_TK[20] WL_TK[21] WL_TK[22] 
+ WL_TK[23] WL_TK[24] WL_TK[25] WL_TK[26] WL_TK[27] WL_TK[28] WL_TK[29] 
+ WL_TK[30] WL_TK[31] NET60[0] NET60[1] NET60[2] NET60[3] NET60[4] NET60[5] 
+ NET60[6] NET60[7] NET59 NET69 NET57[0] NET57[1] NET57[2] NET57[3] NET57[4] 
+ NET57[5] NET57[6] NET57[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
XTRKNORX16_DUMY1 BL_TK VDDI VSSI WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] 
+ WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] 
+ WL_TK[32] WL_TK[33] WL_TK[34] WL_TK[35] WL_TK[36] WL_TK[37] WL_TK[38] 
+ WL_TK[39] WL_TK[40] WL_TK[41] WL_TK[42] WL_TK[43] WL_TK[44] WL_TK[45] 
+ WL_TK[46] WL_TK[47] NET50[0] NET50[1] NET50[2] NET50[3] NET50[4] NET50[5] 
+ NET50[6] NET50[7] NET49 NET59 NET47[0] NET47[1] NET47[2] NET47[3] NET47[4] 
+ NET47[5] NET47[6] NET47[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
XTRKNORX16_BCELL BL_TK VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] 
+ WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL_TK[0] 
+ WL_TK[1] WL_TK[2] WL_TK[3] WL_TK[4] WL_TK[5] WL_TK[6] WL_TK[7] WL_TK[8] 
+ WL_TK[9] WL_TK[10] WL_TK[11] WL_TK[12] WL_TK[13] WL_TK[14] WL_TK[15] 
+ NET70[0] NET70[1] NET70[2] NET70[3] NET70[4] NET70[5] NET70[6] NET70[7] 
+ NET69 NET68 NET67[0] NET67[1] NET67[2] NET67[3] NET67[4] NET67[5] NET67[6] 
+ NET67[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
XTRKNORX16_DUMY2 BL_TK VDDI VSSI WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] 
+ WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] 
+ WL_TK[48] WL_TK[49] WL_TK[50] WL_TK[51] WL_TK[52] WL_TK[53] WL_TK[54] 
+ WL_TK[55] WL_TK[56] WL_TK[57] WL_TK[58] WL_TK[59] WL_TK[60] WL_TK[61] 
+ WL_TK[62] WL_TK[63] NET40[0] NET40[1] NET40[2] NET40[3] NET40[4] NET40[5] 
+ NET40[6] NET40[7] NET39 NET49 NET37[0] NET37[1] NET37[2] NET37[3] NET37[4] 
+ NET37[5] NET37[6] NET37[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    TKBL_S256_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TKBL_S256_CHAR BL_TK VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL_TK[0] 
+ WL_TK[1] WL_TK[2] WL_TK[3] WL_TK[4] WL_TK[5] WL_TK[6] WL_TK[7] WL_TK[8] 
+ WL_TK[9] WL_TK[10] WL_TK[11] WL_TK[12] WL_TK[13] WL_TK[14] WL_TK[15] 
+ WL_TK[16] WL_TK[17] WL_TK[18] WL_TK[19] WL_TK[20] WL_TK[21] WL_TK[22] 
+ WL_TK[23] WL_TK[24] WL_TK[25] WL_TK[26] WL_TK[27] WL_TK[28] WL_TK[29] 
+ WL_TK[30] WL_TK[31] WL_TK[32] WL_TK[33] WL_TK[34] WL_TK[35] WL_TK[36] 
+ WL_TK[37] WL_TK[38] WL_TK[39] WL_TK[40] WL_TK[41] WL_TK[42] WL_TK[43] 
+ WL_TK[44] WL_TK[45] WL_TK[46] WL_TK[47] WL_TK[48] WL_TK[49] WL_TK[50] 
+ WL_TK[51] WL_TK[52] WL_TK[53] WL_TK[54] WL_TK[55] WL_TK[56] WL_TK[57] 
+ WL_TK[58] WL_TK[59] WL_TK[60] WL_TK[61] WL_TK[62] WL_TK[63] WL_TK[64] 
+ WL_TK[65] WL_TK[66] WL_TK[67] WL_TK[68] WL_TK[69] WL_TK[70] WL_TK[71] 
+ WL_TK[72] WL_TK[73] WL_TK[74] WL_TK[75] WL_TK[76] WL_TK[77] WL_TK[78] 
+ WL_TK[79] WL_TK[80] WL_TK[81] WL_TK[82] WL_TK[83] WL_TK[84] WL_TK[85] 
+ WL_TK[86] WL_TK[87] WL_TK[88] WL_TK[89] WL_TK[90] WL_TK[91] WL_TK[92] 
+ WL_TK[93] WL_TK[94] WL_TK[95] WL_TK[96] WL_TK[97] WL_TK[98] WL_TK[99] 
+ WL_TK[100] WL_TK[101] WL_TK[102] WL_TK[103] WL_TK[104] WL_TK[105] WL_TK[106] 
+ WL_TK[107] WL_TK[108] WL_TK[109] WL_TK[110] WL_TK[111] WL_TK[112] WL_TK[113] 
+ WL_TK[114] WL_TK[115] WL_TK[116] WL_TK[117] WL_TK[118] WL_TK[119] WL_TK[120] 
+ WL_TK[121] WL_TK[122] WL_TK[123] WL_TK[124] WL_TK[125] WL_TK[126] WL_TK[127] 
+ WL_TK[128] WL_TK[129] WL_TK[130] WL_TK[131] WL_TK[132] WL_TK[133] WL_TK[134] 
+ WL_TK[135] WL_TK[136] WL_TK[137] WL_TK[138] WL_TK[139] WL_TK[140] WL_TK[141] 
+ WL_TK[142] WL_TK[143] WL_TK[144] WL_TK[145] WL_TK[146] WL_TK[147] WL_TK[148] 
+ WL_TK[149] WL_TK[150] WL_TK[151] WL_TK[152] WL_TK[153] WL_TK[154] WL_TK[155] 
+ WL_TK[156] WL_TK[157] WL_TK[158] WL_TK[159] WL_TK[160] WL_TK[161] WL_TK[162] 
+ WL_TK[163] WL_TK[164] WL_TK[165] WL_TK[166] WL_TK[167] WL_TK[168] WL_TK[169] 
+ WL_TK[170] WL_TK[171] WL_TK[172] WL_TK[173] WL_TK[174] WL_TK[175] WL_TK[176] 
+ WL_TK[177] WL_TK[178] WL_TK[179] WL_TK[180] WL_TK[181] WL_TK[182] WL_TK[183] 
+ WL_TK[184] WL_TK[185] WL_TK[186] WL_TK[187] WL_TK[188] WL_TK[189] WL_TK[190] 
+ WL_TK[191] WL_TK[192] WL_TK[193] WL_TK[194] WL_TK[195] WL_TK[196] WL_TK[197] 
+ WL_TK[198] WL_TK[199] WL_TK[200] WL_TK[201] WL_TK[202] WL_TK[203] WL_TK[204] 
+ WL_TK[205] WL_TK[206] WL_TK[207] WL_TK[208] WL_TK[209] WL_TK[210] WL_TK[211] 
+ WL_TK[212] WL_TK[213] WL_TK[214] WL_TK[215] WL_TK[216] WL_TK[217] WL_TK[218] 
+ WL_TK[219] WL_TK[220] WL_TK[221] WL_TK[222] WL_TK[223] WL_TK[224] WL_TK[225] 
+ WL_TK[226] WL_TK[227] WL_TK[228] WL_TK[229] WL_TK[230] WL_TK[231] WL_TK[232] 
+ WL_TK[233] WL_TK[234] WL_TK[235] WL_TK[236] WL_TK[237] WL_TK[238] WL_TK[239] 
+ WL_TK[240] WL_TK[241] WL_TK[242] WL_TK[243] WL_TK[244] WL_TK[245] WL_TK[246] 
+ WL_TK[247] WL_TK[248] WL_TK[249] WL_TK[250] WL_TK[251] WL_TK[252] WL_TK[253] 
+ WL_TK[254] WL_TK[255] TIEH TIEL
*.PININFO BL_TK:B VDDI:B VSSI:B WL[0]:B WL[1]:B WL[2]:B WL[3]:B WL[4]:B 
*.PININFO WL[5]:B WL[6]:B WL[7]:B WL[8]:B WL[9]:B WL[10]:B WL[11]:B WL[12]:B 
*.PININFO WL[13]:B WL[14]:B WL[15]:B WL[16]:B WL[17]:B WL[18]:B WL[19]:B 
*.PININFO WL[20]:B WL[21]:B WL[22]:B WL[23]:B WL[24]:B WL[25]:B WL[26]:B 
*.PININFO WL[27]:B WL[28]:B WL[29]:B WL[30]:B WL[31]:B WL[32]:B WL[33]:B 
*.PININFO WL[34]:B WL[35]:B WL[36]:B WL[37]:B WL[38]:B WL[39]:B WL[40]:B 
*.PININFO WL[41]:B WL[42]:B WL[43]:B WL[44]:B WL[45]:B WL[46]:B WL[47]:B 
*.PININFO WL[48]:B WL[49]:B WL[50]:B WL[51]:B WL[52]:B WL[53]:B WL[54]:B 
*.PININFO WL[55]:B WL[56]:B WL[57]:B WL[58]:B WL[59]:B WL[60]:B WL[61]:B 
*.PININFO WL[62]:B WL[63]:B WL[64]:B WL[65]:B WL[66]:B WL[67]:B WL[68]:B 
*.PININFO WL[69]:B WL[70]:B WL[71]:B WL[72]:B WL[73]:B WL[74]:B WL[75]:B 
*.PININFO WL[76]:B WL[77]:B WL[78]:B WL[79]:B WL[80]:B WL[81]:B WL[82]:B 
*.PININFO WL[83]:B WL[84]:B WL[85]:B WL[86]:B WL[87]:B WL[88]:B WL[89]:B 
*.PININFO WL[90]:B WL[91]:B WL[92]:B WL[93]:B WL[94]:B WL[95]:B WL[96]:B 
*.PININFO WL[97]:B WL[98]:B WL[99]:B WL[100]:B WL[101]:B WL[102]:B WL[103]:B 
*.PININFO WL[104]:B WL[105]:B WL[106]:B WL[107]:B WL[108]:B WL[109]:B 
*.PININFO WL[110]:B WL[111]:B WL[112]:B WL[113]:B WL[114]:B WL[115]:B 
*.PININFO WL[116]:B WL[117]:B WL[118]:B WL[119]:B WL[120]:B WL[121]:B 
*.PININFO WL[122]:B WL[123]:B WL[124]:B WL[125]:B WL[126]:B WL[127]:B 
*.PININFO WL[128]:B WL[129]:B WL[130]:B WL[131]:B WL[132]:B WL[133]:B 
*.PININFO WL[134]:B WL[135]:B WL[136]:B WL[137]:B WL[138]:B WL[139]:B 
*.PININFO WL[140]:B WL[141]:B WL[142]:B WL[143]:B WL[144]:B WL[145]:B 
*.PININFO WL[146]:B WL[147]:B WL[148]:B WL[149]:B WL[150]:B WL[151]:B 
*.PININFO WL[152]:B WL[153]:B WL[154]:B WL[155]:B WL[156]:B WL[157]:B 
*.PININFO WL[158]:B WL[159]:B WL[160]:B WL[161]:B WL[162]:B WL[163]:B 
*.PININFO WL[164]:B WL[165]:B WL[166]:B WL[167]:B WL[168]:B WL[169]:B 
*.PININFO WL[170]:B WL[171]:B WL[172]:B WL[173]:B WL[174]:B WL[175]:B 
*.PININFO WL[176]:B WL[177]:B WL[178]:B WL[179]:B WL[180]:B WL[181]:B 
*.PININFO WL[182]:B WL[183]:B WL[184]:B WL[185]:B WL[186]:B WL[187]:B 
*.PININFO WL[188]:B WL[189]:B WL[190]:B WL[191]:B WL[192]:B WL[193]:B 
*.PININFO WL[194]:B WL[195]:B WL[196]:B WL[197]:B WL[198]:B WL[199]:B 
*.PININFO WL[200]:B WL[201]:B WL[202]:B WL[203]:B WL[204]:B WL[205]:B 
*.PININFO WL[206]:B WL[207]:B WL[208]:B WL[209]:B WL[210]:B WL[211]:B 
*.PININFO WL[212]:B WL[213]:B WL[214]:B WL[215]:B WL[216]:B WL[217]:B 
*.PININFO WL[218]:B WL[219]:B WL[220]:B WL[221]:B WL[222]:B WL[223]:B 
*.PININFO WL[224]:B WL[225]:B WL[226]:B WL[227]:B WL[228]:B WL[229]:B 
*.PININFO WL[230]:B WL[231]:B WL[232]:B WL[233]:B WL[234]:B WL[235]:B 
*.PININFO WL[236]:B WL[237]:B WL[238]:B WL[239]:B WL[240]:B WL[241]:B 
*.PININFO WL[242]:B WL[243]:B WL[244]:B WL[245]:B WL[246]:B WL[247]:B 
*.PININFO WL[248]:B WL[249]:B WL[250]:B WL[251]:B WL[252]:B WL[253]:B 
*.PININFO WL[254]:B WL[255]:B WL_TK[0]:B WL_TK[1]:B WL_TK[2]:B WL_TK[3]:B 
*.PININFO WL_TK[4]:B WL_TK[5]:B WL_TK[6]:B WL_TK[7]:B WL_TK[8]:B WL_TK[9]:B 
*.PININFO WL_TK[10]:B WL_TK[11]:B WL_TK[12]:B WL_TK[13]:B WL_TK[14]:B 
*.PININFO WL_TK[15]:B WL_TK[16]:B WL_TK[17]:B WL_TK[18]:B WL_TK[19]:B 
*.PININFO WL_TK[20]:B WL_TK[21]:B WL_TK[22]:B WL_TK[23]:B WL_TK[24]:B 
*.PININFO WL_TK[25]:B WL_TK[26]:B WL_TK[27]:B WL_TK[28]:B WL_TK[29]:B 
*.PININFO WL_TK[30]:B WL_TK[31]:B WL_TK[32]:B WL_TK[33]:B WL_TK[34]:B 
*.PININFO WL_TK[35]:B WL_TK[36]:B WL_TK[37]:B WL_TK[38]:B WL_TK[39]:B 
*.PININFO WL_TK[40]:B WL_TK[41]:B WL_TK[42]:B WL_TK[43]:B WL_TK[44]:B 
*.PININFO WL_TK[45]:B WL_TK[46]:B WL_TK[47]:B WL_TK[48]:B WL_TK[49]:B 
*.PININFO WL_TK[50]:B WL_TK[51]:B WL_TK[52]:B WL_TK[53]:B WL_TK[54]:B 
*.PININFO WL_TK[55]:B WL_TK[56]:B WL_TK[57]:B WL_TK[58]:B WL_TK[59]:B 
*.PININFO WL_TK[60]:B WL_TK[61]:B WL_TK[62]:B WL_TK[63]:B WL_TK[64]:B 
*.PININFO WL_TK[65]:B WL_TK[66]:B WL_TK[67]:B WL_TK[68]:B WL_TK[69]:B 
*.PININFO WL_TK[70]:B WL_TK[71]:B WL_TK[72]:B WL_TK[73]:B WL_TK[74]:B 
*.PININFO WL_TK[75]:B WL_TK[76]:B WL_TK[77]:B WL_TK[78]:B WL_TK[79]:B 
*.PININFO WL_TK[80]:B WL_TK[81]:B WL_TK[82]:B WL_TK[83]:B WL_TK[84]:B 
*.PININFO WL_TK[85]:B WL_TK[86]:B WL_TK[87]:B WL_TK[88]:B WL_TK[89]:B 
*.PININFO WL_TK[90]:B WL_TK[91]:B WL_TK[92]:B WL_TK[93]:B WL_TK[94]:B 
*.PININFO WL_TK[95]:B WL_TK[96]:B WL_TK[97]:B WL_TK[98]:B WL_TK[99]:B 
*.PININFO WL_TK[100]:B WL_TK[101]:B WL_TK[102]:B WL_TK[103]:B WL_TK[104]:B 
*.PININFO WL_TK[105]:B WL_TK[106]:B WL_TK[107]:B WL_TK[108]:B WL_TK[109]:B 
*.PININFO WL_TK[110]:B WL_TK[111]:B WL_TK[112]:B WL_TK[113]:B WL_TK[114]:B 
*.PININFO WL_TK[115]:B WL_TK[116]:B WL_TK[117]:B WL_TK[118]:B WL_TK[119]:B 
*.PININFO WL_TK[120]:B WL_TK[121]:B WL_TK[122]:B WL_TK[123]:B WL_TK[124]:B 
*.PININFO WL_TK[125]:B WL_TK[126]:B WL_TK[127]:B WL_TK[128]:B WL_TK[129]:B 
*.PININFO WL_TK[130]:B WL_TK[131]:B WL_TK[132]:B WL_TK[133]:B WL_TK[134]:B 
*.PININFO WL_TK[135]:B WL_TK[136]:B WL_TK[137]:B WL_TK[138]:B WL_TK[139]:B 
*.PININFO WL_TK[140]:B WL_TK[141]:B WL_TK[142]:B WL_TK[143]:B WL_TK[144]:B 
*.PININFO WL_TK[145]:B WL_TK[146]:B WL_TK[147]:B WL_TK[148]:B WL_TK[149]:B 
*.PININFO WL_TK[150]:B WL_TK[151]:B WL_TK[152]:B WL_TK[153]:B WL_TK[154]:B 
*.PININFO WL_TK[155]:B WL_TK[156]:B WL_TK[157]:B WL_TK[158]:B WL_TK[159]:B 
*.PININFO WL_TK[160]:B WL_TK[161]:B WL_TK[162]:B WL_TK[163]:B WL_TK[164]:B 
*.PININFO WL_TK[165]:B WL_TK[166]:B WL_TK[167]:B WL_TK[168]:B WL_TK[169]:B 
*.PININFO WL_TK[170]:B WL_TK[171]:B WL_TK[172]:B WL_TK[173]:B WL_TK[174]:B 
*.PININFO WL_TK[175]:B WL_TK[176]:B WL_TK[177]:B WL_TK[178]:B WL_TK[179]:B 
*.PININFO WL_TK[180]:B WL_TK[181]:B WL_TK[182]:B WL_TK[183]:B WL_TK[184]:B 
*.PININFO WL_TK[185]:B WL_TK[186]:B WL_TK[187]:B WL_TK[188]:B WL_TK[189]:B 
*.PININFO WL_TK[190]:B WL_TK[191]:B WL_TK[192]:B WL_TK[193]:B WL_TK[194]:B 
*.PININFO WL_TK[195]:B WL_TK[196]:B WL_TK[197]:B WL_TK[198]:B WL_TK[199]:B 
*.PININFO WL_TK[200]:B WL_TK[201]:B WL_TK[202]:B WL_TK[203]:B WL_TK[204]:B 
*.PININFO WL_TK[205]:B WL_TK[206]:B WL_TK[207]:B WL_TK[208]:B WL_TK[209]:B 
*.PININFO WL_TK[210]:B WL_TK[211]:B WL_TK[212]:B WL_TK[213]:B WL_TK[214]:B 
*.PININFO WL_TK[215]:B WL_TK[216]:B WL_TK[217]:B WL_TK[218]:B WL_TK[219]:B 
*.PININFO WL_TK[220]:B WL_TK[221]:B WL_TK[222]:B WL_TK[223]:B WL_TK[224]:B 
*.PININFO WL_TK[225]:B WL_TK[226]:B WL_TK[227]:B WL_TK[228]:B WL_TK[229]:B 
*.PININFO WL_TK[230]:B WL_TK[231]:B WL_TK[232]:B WL_TK[233]:B WL_TK[234]:B 
*.PININFO WL_TK[235]:B WL_TK[236]:B WL_TK[237]:B WL_TK[238]:B WL_TK[239]:B 
*.PININFO WL_TK[240]:B WL_TK[241]:B WL_TK[242]:B WL_TK[243]:B WL_TK[244]:B 
*.PININFO WL_TK[245]:B WL_TK[246]:B WL_TK[247]:B WL_TK[248]:B WL_TK[249]:B 
*.PININFO WL_TK[250]:B WL_TK[251]:B WL_TK[252]:B WL_TK[253]:B WL_TK[254]:B 
*.PININFO WL_TK[255]:B TIEH:B TIEL:B
XTRKNORX64_DUMY4 BL_TK VDDI VSSI WL[128] WL[129] WL[130] WL[131] WL[132] 
+ WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] WL[140] WL[141] 
+ WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] WL[149] WL[150] 
+ WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] WL[158] WL[159] 
+ WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] WL[167] WL[168] 
+ WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] WL[176] WL[177] 
+ WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] WL[185] WL[186] 
+ WL[187] WL[188] WL[189] WL[190] WL[191] WL_TK[128] WL_TK[129] WL_TK[130] 
+ WL_TK[131] WL_TK[132] WL_TK[133] WL_TK[134] WL_TK[135] WL_TK[136] WL_TK[137] 
+ WL_TK[138] WL_TK[139] WL_TK[140] WL_TK[141] WL_TK[142] WL_TK[143] WL_TK[144] 
+ WL_TK[145] WL_TK[146] WL_TK[147] WL_TK[148] WL_TK[149] WL_TK[150] WL_TK[151] 
+ WL_TK[152] WL_TK[153] WL_TK[154] WL_TK[155] WL_TK[156] WL_TK[157] WL_TK[158] 
+ WL_TK[159] WL_TK[160] WL_TK[161] WL_TK[162] WL_TK[163] WL_TK[164] WL_TK[165] 
+ WL_TK[166] WL_TK[167] WL_TK[168] WL_TK[169] WL_TK[170] WL_TK[171] WL_TK[172] 
+ WL_TK[173] WL_TK[174] WL_TK[175] WL_TK[176] WL_TK[177] WL_TK[178] WL_TK[179] 
+ WL_TK[180] WL_TK[181] WL_TK[182] WL_TK[183] WL_TK[184] WL_TK[185] WL_TK[186] 
+ WL_TK[187] WL_TK[188] WL_TK[189] WL_TK[190] WL_TK[191] NET20[0] NET20[1] 
+ NET20[2] NET20[3] NET20[4] NET20[5] NET20[6] NET20[7] NET20[8] NET20[9] 
+ NET20[10] NET20[11] NET20[12] NET20[13] NET20[14] NET20[15] NET20[16] 
+ NET20[17] NET20[18] NET20[19] NET20[20] NET20[21] NET20[22] NET20[23] 
+ NET20[24] NET20[25] NET20[26] NET20[27] NET20[28] NET20[29] NET20[30] 
+ NET20[31] NET19 NET18 NET17[0] NET17[1] NET17[2] NET17[3] NET17[4] NET17[5] 
+ NET17[6] NET17[7] NET17[8] NET17[9] NET17[10] NET17[11] NET17[12] NET17[13] 
+ NET17[14] NET17[15] NET17[16] NET17[17] NET17[18] NET17[19] NET17[20] 
+ NET17[21] NET17[22] NET17[23] NET17[24] NET17[25] NET17[26] NET17[27] 
+ NET17[28] NET17[29] NET17[30] NET17[31] TIEH S1AHSF400W40_TRKNORX64_CHAR
XTRKNORX64_DUMY3 BL_TK VDDI VSSI WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] 
+ WL[70] WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] 
+ WL[81] WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] 
+ WL[92] WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] 
+ WL[102] WL[103] WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] 
+ WL[111] WL[112] WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] 
+ WL[120] WL[121] WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL_TK[64] 
+ WL_TK[65] WL_TK[66] WL_TK[67] WL_TK[68] WL_TK[69] WL_TK[70] WL_TK[71] 
+ WL_TK[72] WL_TK[73] WL_TK[74] WL_TK[75] WL_TK[76] WL_TK[77] WL_TK[78] 
+ WL_TK[79] WL_TK[80] WL_TK[81] WL_TK[82] WL_TK[83] WL_TK[84] WL_TK[85] 
+ WL_TK[86] WL_TK[87] WL_TK[88] WL_TK[89] WL_TK[90] WL_TK[91] WL_TK[92] 
+ WL_TK[93] WL_TK[94] WL_TK[95] WL_TK[96] WL_TK[97] WL_TK[98] WL_TK[99] 
+ WL_TK[100] WL_TK[101] WL_TK[102] WL_TK[103] WL_TK[104] WL_TK[105] WL_TK[106] 
+ WL_TK[107] WL_TK[108] WL_TK[109] WL_TK[110] WL_TK[111] WL_TK[112] WL_TK[113] 
+ WL_TK[114] WL_TK[115] WL_TK[116] WL_TK[117] WL_TK[118] WL_TK[119] WL_TK[120] 
+ WL_TK[121] WL_TK[122] WL_TK[123] WL_TK[124] WL_TK[125] WL_TK[126] WL_TK[127] 
+ NET10[0] NET10[1] NET10[2] NET10[3] NET10[4] NET10[5] NET10[6] NET10[7] 
+ NET10[8] NET10[9] NET10[10] NET10[11] NET10[12] NET10[13] NET10[14] 
+ NET10[15] NET10[16] NET10[17] NET10[18] NET10[19] NET10[20] NET10[21] 
+ NET10[22] NET10[23] NET10[24] NET10[25] NET10[26] NET10[27] NET10[28] 
+ NET10[29] NET10[30] NET10[31] NET9 NET8 NET7[0] NET7[1] NET7[2] NET7[3] 
+ NET7[4] NET7[5] NET7[6] NET7[7] NET7[8] NET7[9] NET7[10] NET7[11] NET7[12] 
+ NET7[13] NET7[14] NET7[15] NET7[16] NET7[17] NET7[18] NET7[19] NET7[20] 
+ NET7[21] NET7[22] NET7[23] NET7[24] NET7[25] NET7[26] NET7[27] NET7[28] 
+ NET7[29] NET7[30] NET7[31] TIEH S1AHSF400W40_TRKNORX64_CHAR
XTRKNORX64_DYMY5 BL_TK VDDI VSSI WL[192] WL[193] WL[194] WL[195] WL[196] 
+ WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] WL[203] WL[204] WL[205] 
+ WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] WL[212] WL[213] WL[214] 
+ WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] WL[221] WL[222] WL[223] 
+ WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] WL[230] WL[231] WL[232] 
+ WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] WL[239] WL[240] WL[241] 
+ WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] WL[248] WL[249] WL[250] 
+ WL[251] WL[252] WL[253] WL[254] WL[255] WL_TK[192] WL_TK[193] WL_TK[194] 
+ WL_TK[195] WL_TK[196] WL_TK[197] WL_TK[198] WL_TK[199] WL_TK[200] WL_TK[201] 
+ WL_TK[202] WL_TK[203] WL_TK[204] WL_TK[205] WL_TK[206] WL_TK[207] WL_TK[208] 
+ WL_TK[209] WL_TK[210] WL_TK[211] WL_TK[212] WL_TK[213] WL_TK[214] WL_TK[215] 
+ WL_TK[216] WL_TK[217] WL_TK[218] WL_TK[219] WL_TK[220] WL_TK[221] WL_TK[222] 
+ WL_TK[223] WL_TK[224] WL_TK[225] WL_TK[226] WL_TK[227] WL_TK[228] WL_TK[229] 
+ WL_TK[230] WL_TK[231] WL_TK[232] WL_TK[233] WL_TK[234] WL_TK[235] WL_TK[236] 
+ WL_TK[237] WL_TK[238] WL_TK[239] WL_TK[240] WL_TK[241] WL_TK[242] WL_TK[243] 
+ WL_TK[244] WL_TK[245] WL_TK[246] WL_TK[247] WL_TK[248] WL_TK[249] WL_TK[250] 
+ WL_TK[251] WL_TK[252] WL_TK[253] WL_TK[254] WL_TK[255] NET30[0] NET30[1] 
+ NET30[2] NET30[3] NET30[4] NET30[5] NET30[6] NET30[7] NET30[8] NET30[9] 
+ NET30[10] NET30[11] NET30[12] NET30[13] NET30[14] NET30[15] NET30[16] 
+ NET30[17] NET30[18] NET30[19] NET30[20] NET30[21] NET30[22] NET30[23] 
+ NET30[24] NET30[25] NET30[26] NET30[27] NET30[28] NET30[29] NET30[30] 
+ NET30[31] NET29 NET28 NET27[0] NET27[1] NET27[2] NET27[3] NET27[4] NET27[5] 
+ NET27[6] NET27[7] NET27[8] NET27[9] NET27[10] NET27[11] NET27[12] NET27[13] 
+ NET27[14] NET27[15] NET27[16] NET27[17] NET27[18] NET27[19] NET27[20] 
+ NET27[21] NET27[22] NET27[23] NET27[24] NET27[25] NET27[26] NET27[27] 
+ NET27[28] NET27[29] NET27[30] NET27[31] TIEH S1AHSF400W40_TRKNORX64_CHAR
XTRKNORX16_DUMY0 BL_TK VDDI VSSI WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] 
+ WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] 
+ WL_TK[16] WL_TK[17] WL_TK[18] WL_TK[19] WL_TK[20] WL_TK[21] WL_TK[22] 
+ WL_TK[23] WL_TK[24] WL_TK[25] WL_TK[26] WL_TK[27] WL_TK[28] WL_TK[29] 
+ WL_TK[30] WL_TK[31] NET60[0] NET60[1] NET60[2] NET60[3] NET60[4] NET60[5] 
+ NET60[6] NET60[7] NET59 NET69 NET57[0] NET57[1] NET57[2] NET57[3] NET57[4] 
+ NET57[5] NET57[6] NET57[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
XTRKNORX16_DUMY1 BL_TK VDDI VSSI WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] 
+ WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] 
+ WL_TK[32] WL_TK[33] WL_TK[34] WL_TK[35] WL_TK[36] WL_TK[37] WL_TK[38] 
+ WL_TK[39] WL_TK[40] WL_TK[41] WL_TK[42] WL_TK[43] WL_TK[44] WL_TK[45] 
+ WL_TK[46] WL_TK[47] NET50[0] NET50[1] NET50[2] NET50[3] NET50[4] NET50[5] 
+ NET50[6] NET50[7] NET49 NET59 NET47[0] NET47[1] NET47[2] NET47[3] NET47[4] 
+ NET47[5] NET47[6] NET47[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
XTRKNORX16_BCELL BL_TK VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] 
+ WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL_TK[0] 
+ WL_TK[1] WL_TK[2] WL_TK[3] WL_TK[4] WL_TK[5] WL_TK[6] WL_TK[7] WL_TK[8] 
+ WL_TK[9] WL_TK[10] WL_TK[11] WL_TK[12] WL_TK[13] WL_TK[14] WL_TK[15] 
+ NET70[0] NET70[1] NET70[2] NET70[3] NET70[4] NET70[5] NET70[6] NET70[7] 
+ NET69 NET68 NET67[0] NET67[1] NET67[2] NET67[3] NET67[4] NET67[5] NET67[6] 
+ NET67[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
XTRKNORX16_DUMY2 BL_TK VDDI VSSI WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] 
+ WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] 
+ WL_TK[48] WL_TK[49] WL_TK[50] WL_TK[51] WL_TK[52] WL_TK[53] WL_TK[54] 
+ WL_TK[55] WL_TK[56] WL_TK[57] WL_TK[58] WL_TK[59] WL_TK[60] WL_TK[61] 
+ WL_TK[62] WL_TK[63] NET40[0] NET40[1] NET40[2] NET40[3] NET40[4] NET40[5] 
+ NET40[6] NET40[7] NET39 NET49 NET37[0] NET37[1] NET37[2] NET37[3] NET37[4] 
+ NET37[5] NET37[6] NET37[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    TKBL_S32_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TKBL_S32_CHAR BL_TK VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL_TK[0] WL_TK[1] WL_TK[2] WL_TK[3] WL_TK[4] 
+ WL_TK[5] WL_TK[6] WL_TK[7] WL_TK[8] WL_TK[9] WL_TK[10] WL_TK[11] WL_TK[12] 
+ WL_TK[13] WL_TK[14] WL_TK[15] WL_TK[16] WL_TK[17] WL_TK[18] WL_TK[19] 
+ WL_TK[20] WL_TK[21] WL_TK[22] WL_TK[23] WL_TK[24] WL_TK[25] WL_TK[26] 
+ WL_TK[27] WL_TK[28] WL_TK[29] WL_TK[30] WL_TK[31] TIEH TIEL
*.PININFO BL_TK:B VDDI:B VSSI:B WL[0]:B WL[1]:B WL[2]:B WL[3]:B WL[4]:B 
*.PININFO WL[5]:B WL[6]:B WL[7]:B WL[8]:B WL[9]:B WL[10]:B WL[11]:B WL[12]:B 
*.PININFO WL[13]:B WL[14]:B WL[15]:B WL[16]:B WL[17]:B WL[18]:B WL[19]:B 
*.PININFO WL[20]:B WL[21]:B WL[22]:B WL[23]:B WL[24]:B WL[25]:B WL[26]:B 
*.PININFO WL[27]:B WL[28]:B WL[29]:B WL[30]:B WL[31]:B WL_TK[0]:B WL_TK[1]:B 
*.PININFO WL_TK[2]:B WL_TK[3]:B WL_TK[4]:B WL_TK[5]:B WL_TK[6]:B WL_TK[7]:B 
*.PININFO WL_TK[8]:B WL_TK[9]:B WL_TK[10]:B WL_TK[11]:B WL_TK[12]:B 
*.PININFO WL_TK[13]:B WL_TK[14]:B WL_TK[15]:B WL_TK[16]:B WL_TK[17]:B 
*.PININFO WL_TK[18]:B WL_TK[19]:B WL_TK[20]:B WL_TK[21]:B WL_TK[22]:B 
*.PININFO WL_TK[23]:B WL_TK[24]:B WL_TK[25]:B WL_TK[26]:B WL_TK[27]:B 
*.PININFO WL_TK[28]:B WL_TK[29]:B WL_TK[30]:B WL_TK[31]:B TIEH:B TIEL:B
XTRKNORX16_DUMY0 BL_TK VDDI VSSI WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] 
+ WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] 
+ WL_TK[16] WL_TK[17] WL_TK[18] WL_TK[19] WL_TK[20] WL_TK[21] WL_TK[22] 
+ WL_TK[23] WL_TK[24] WL_TK[25] WL_TK[26] WL_TK[27] WL_TK[28] WL_TK[29] 
+ WL_TK[30] WL_TK[31] NET60[0] NET60[1] NET60[2] NET60[3] NET60[4] NET60[5] 
+ NET60[6] NET60[7] NET59 NET69 NET57[0] NET57[1] NET57[2] NET57[3] NET57[4] 
+ NET57[5] NET57[6] NET57[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
XTRKNORX16_BCELL BL_TK VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] 
+ WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL_TK[0] 
+ WL_TK[1] WL_TK[2] WL_TK[3] WL_TK[4] WL_TK[5] WL_TK[6] WL_TK[7] WL_TK[8] 
+ WL_TK[9] WL_TK[10] WL_TK[11] WL_TK[12] WL_TK[13] WL_TK[14] WL_TK[15] 
+ NET70[0] NET70[1] NET70[2] NET70[3] NET70[4] NET70[5] NET70[6] NET70[7] 
+ NET69 NET68 NET67[0] NET67[1] NET67[2] NET67[3] NET67[4] NET67[5] NET67[6] 
+ NET67[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    TKBL_S128_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TKBL_S128_CHAR BL_TK VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL_TK[0] WL_TK[1] WL_TK[2] 
+ WL_TK[3] WL_TK[4] WL_TK[5] WL_TK[6] WL_TK[7] WL_TK[8] WL_TK[9] WL_TK[10] 
+ WL_TK[11] WL_TK[12] WL_TK[13] WL_TK[14] WL_TK[15] WL_TK[16] WL_TK[17] 
+ WL_TK[18] WL_TK[19] WL_TK[20] WL_TK[21] WL_TK[22] WL_TK[23] WL_TK[24] 
+ WL_TK[25] WL_TK[26] WL_TK[27] WL_TK[28] WL_TK[29] WL_TK[30] WL_TK[31] 
+ WL_TK[32] WL_TK[33] WL_TK[34] WL_TK[35] WL_TK[36] WL_TK[37] WL_TK[38] 
+ WL_TK[39] WL_TK[40] WL_TK[41] WL_TK[42] WL_TK[43] WL_TK[44] WL_TK[45] 
+ WL_TK[46] WL_TK[47] WL_TK[48] WL_TK[49] WL_TK[50] WL_TK[51] WL_TK[52] 
+ WL_TK[53] WL_TK[54] WL_TK[55] WL_TK[56] WL_TK[57] WL_TK[58] WL_TK[59] 
+ WL_TK[60] WL_TK[61] WL_TK[62] WL_TK[63] WL_TK[64] WL_TK[65] WL_TK[66] 
+ WL_TK[67] WL_TK[68] WL_TK[69] WL_TK[70] WL_TK[71] WL_TK[72] WL_TK[73] 
+ WL_TK[74] WL_TK[75] WL_TK[76] WL_TK[77] WL_TK[78] WL_TK[79] WL_TK[80] 
+ WL_TK[81] WL_TK[82] WL_TK[83] WL_TK[84] WL_TK[85] WL_TK[86] WL_TK[87] 
+ WL_TK[88] WL_TK[89] WL_TK[90] WL_TK[91] WL_TK[92] WL_TK[93] WL_TK[94] 
+ WL_TK[95] WL_TK[96] WL_TK[97] WL_TK[98] WL_TK[99] WL_TK[100] WL_TK[101] 
+ WL_TK[102] WL_TK[103] WL_TK[104] WL_TK[105] WL_TK[106] WL_TK[107] WL_TK[108] 
+ WL_TK[109] WL_TK[110] WL_TK[111] WL_TK[112] WL_TK[113] WL_TK[114] WL_TK[115] 
+ WL_TK[116] WL_TK[117] WL_TK[118] WL_TK[119] WL_TK[120] WL_TK[121] WL_TK[122] 
+ WL_TK[123] WL_TK[124] WL_TK[125] WL_TK[126] WL_TK[127] TIEH TIEL
*.PININFO BL_TK:B VDDI:B VSSI:B WL[0]:B WL[1]:B WL[2]:B WL[3]:B WL[4]:B 
*.PININFO WL[5]:B WL[6]:B WL[7]:B WL[8]:B WL[9]:B WL[10]:B WL[11]:B WL[12]:B 
*.PININFO WL[13]:B WL[14]:B WL[15]:B WL[16]:B WL[17]:B WL[18]:B WL[19]:B 
*.PININFO WL[20]:B WL[21]:B WL[22]:B WL[23]:B WL[24]:B WL[25]:B WL[26]:B 
*.PININFO WL[27]:B WL[28]:B WL[29]:B WL[30]:B WL[31]:B WL[32]:B WL[33]:B 
*.PININFO WL[34]:B WL[35]:B WL[36]:B WL[37]:B WL[38]:B WL[39]:B WL[40]:B 
*.PININFO WL[41]:B WL[42]:B WL[43]:B WL[44]:B WL[45]:B WL[46]:B WL[47]:B 
*.PININFO WL[48]:B WL[49]:B WL[50]:B WL[51]:B WL[52]:B WL[53]:B WL[54]:B 
*.PININFO WL[55]:B WL[56]:B WL[57]:B WL[58]:B WL[59]:B WL[60]:B WL[61]:B 
*.PININFO WL[62]:B WL[63]:B WL[64]:B WL[65]:B WL[66]:B WL[67]:B WL[68]:B 
*.PININFO WL[69]:B WL[70]:B WL[71]:B WL[72]:B WL[73]:B WL[74]:B WL[75]:B 
*.PININFO WL[76]:B WL[77]:B WL[78]:B WL[79]:B WL[80]:B WL[81]:B WL[82]:B 
*.PININFO WL[83]:B WL[84]:B WL[85]:B WL[86]:B WL[87]:B WL[88]:B WL[89]:B 
*.PININFO WL[90]:B WL[91]:B WL[92]:B WL[93]:B WL[94]:B WL[95]:B WL[96]:B 
*.PININFO WL[97]:B WL[98]:B WL[99]:B WL[100]:B WL[101]:B WL[102]:B WL[103]:B 
*.PININFO WL[104]:B WL[105]:B WL[106]:B WL[107]:B WL[108]:B WL[109]:B 
*.PININFO WL[110]:B WL[111]:B WL[112]:B WL[113]:B WL[114]:B WL[115]:B 
*.PININFO WL[116]:B WL[117]:B WL[118]:B WL[119]:B WL[120]:B WL[121]:B 
*.PININFO WL[122]:B WL[123]:B WL[124]:B WL[125]:B WL[126]:B WL[127]:B 
*.PININFO WL_TK[0]:B WL_TK[1]:B WL_TK[2]:B WL_TK[3]:B WL_TK[4]:B WL_TK[5]:B 
*.PININFO WL_TK[6]:B WL_TK[7]:B WL_TK[8]:B WL_TK[9]:B WL_TK[10]:B WL_TK[11]:B 
*.PININFO WL_TK[12]:B WL_TK[13]:B WL_TK[14]:B WL_TK[15]:B WL_TK[16]:B 
*.PININFO WL_TK[17]:B WL_TK[18]:B WL_TK[19]:B WL_TK[20]:B WL_TK[21]:B 
*.PININFO WL_TK[22]:B WL_TK[23]:B WL_TK[24]:B WL_TK[25]:B WL_TK[26]:B 
*.PININFO WL_TK[27]:B WL_TK[28]:B WL_TK[29]:B WL_TK[30]:B WL_TK[31]:B 
*.PININFO WL_TK[32]:B WL_TK[33]:B WL_TK[34]:B WL_TK[35]:B WL_TK[36]:B 
*.PININFO WL_TK[37]:B WL_TK[38]:B WL_TK[39]:B WL_TK[40]:B WL_TK[41]:B 
*.PININFO WL_TK[42]:B WL_TK[43]:B WL_TK[44]:B WL_TK[45]:B WL_TK[46]:B 
*.PININFO WL_TK[47]:B WL_TK[48]:B WL_TK[49]:B WL_TK[50]:B WL_TK[51]:B 
*.PININFO WL_TK[52]:B WL_TK[53]:B WL_TK[54]:B WL_TK[55]:B WL_TK[56]:B 
*.PININFO WL_TK[57]:B WL_TK[58]:B WL_TK[59]:B WL_TK[60]:B WL_TK[61]:B 
*.PININFO WL_TK[62]:B WL_TK[63]:B WL_TK[64]:B WL_TK[65]:B WL_TK[66]:B 
*.PININFO WL_TK[67]:B WL_TK[68]:B WL_TK[69]:B WL_TK[70]:B WL_TK[71]:B 
*.PININFO WL_TK[72]:B WL_TK[73]:B WL_TK[74]:B WL_TK[75]:B WL_TK[76]:B 
*.PININFO WL_TK[77]:B WL_TK[78]:B WL_TK[79]:B WL_TK[80]:B WL_TK[81]:B 
*.PININFO WL_TK[82]:B WL_TK[83]:B WL_TK[84]:B WL_TK[85]:B WL_TK[86]:B 
*.PININFO WL_TK[87]:B WL_TK[88]:B WL_TK[89]:B WL_TK[90]:B WL_TK[91]:B 
*.PININFO WL_TK[92]:B WL_TK[93]:B WL_TK[94]:B WL_TK[95]:B WL_TK[96]:B 
*.PININFO WL_TK[97]:B WL_TK[98]:B WL_TK[99]:B WL_TK[100]:B WL_TK[101]:B 
*.PININFO WL_TK[102]:B WL_TK[103]:B WL_TK[104]:B WL_TK[105]:B WL_TK[106]:B 
*.PININFO WL_TK[107]:B WL_TK[108]:B WL_TK[109]:B WL_TK[110]:B WL_TK[111]:B 
*.PININFO WL_TK[112]:B WL_TK[113]:B WL_TK[114]:B WL_TK[115]:B WL_TK[116]:B 
*.PININFO WL_TK[117]:B WL_TK[118]:B WL_TK[119]:B WL_TK[120]:B WL_TK[121]:B 
*.PININFO WL_TK[122]:B WL_TK[123]:B WL_TK[124]:B WL_TK[125]:B WL_TK[126]:B 
*.PININFO WL_TK[127]:B TIEH:B TIEL:B
XTRKNORX64_DUMY3 BL_TK VDDI VSSI WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] 
+ WL[70] WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] 
+ WL[81] WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] 
+ WL[92] WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] 
+ WL[102] WL[103] WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] 
+ WL[111] WL[112] WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] 
+ WL[120] WL[121] WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL_TK[64] 
+ WL_TK[65] WL_TK[66] WL_TK[67] WL_TK[68] WL_TK[69] WL_TK[70] WL_TK[71] 
+ WL_TK[72] WL_TK[73] WL_TK[74] WL_TK[75] WL_TK[76] WL_TK[77] WL_TK[78] 
+ WL_TK[79] WL_TK[80] WL_TK[81] WL_TK[82] WL_TK[83] WL_TK[84] WL_TK[85] 
+ WL_TK[86] WL_TK[87] WL_TK[88] WL_TK[89] WL_TK[90] WL_TK[91] WL_TK[92] 
+ WL_TK[93] WL_TK[94] WL_TK[95] WL_TK[96] WL_TK[97] WL_TK[98] WL_TK[99] 
+ WL_TK[100] WL_TK[101] WL_TK[102] WL_TK[103] WL_TK[104] WL_TK[105] WL_TK[106] 
+ WL_TK[107] WL_TK[108] WL_TK[109] WL_TK[110] WL_TK[111] WL_TK[112] WL_TK[113] 
+ WL_TK[114] WL_TK[115] WL_TK[116] WL_TK[117] WL_TK[118] WL_TK[119] WL_TK[120] 
+ WL_TK[121] WL_TK[122] WL_TK[123] WL_TK[124] WL_TK[125] WL_TK[126] WL_TK[127] 
+ NET10[0] NET10[1] NET10[2] NET10[3] NET10[4] NET10[5] NET10[6] NET10[7] 
+ NET10[8] NET10[9] NET10[10] NET10[11] NET10[12] NET10[13] NET10[14] 
+ NET10[15] NET10[16] NET10[17] NET10[18] NET10[19] NET10[20] NET10[21] 
+ NET10[22] NET10[23] NET10[24] NET10[25] NET10[26] NET10[27] NET10[28] 
+ NET10[29] NET10[30] NET10[31] NET9 NET8 NET7[0] NET7[1] NET7[2] NET7[3] 
+ NET7[4] NET7[5] NET7[6] NET7[7] NET7[8] NET7[9] NET7[10] NET7[11] NET7[12] 
+ NET7[13] NET7[14] NET7[15] NET7[16] NET7[17] NET7[18] NET7[19] NET7[20] 
+ NET7[21] NET7[22] NET7[23] NET7[24] NET7[25] NET7[26] NET7[27] NET7[28] 
+ NET7[29] NET7[30] NET7[31] TIEH S1AHSF400W40_TRKNORX64_CHAR
XTRKNORX16_DUMY0 BL_TK VDDI VSSI WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] 
+ WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] 
+ WL_TK[16] WL_TK[17] WL_TK[18] WL_TK[19] WL_TK[20] WL_TK[21] WL_TK[22] 
+ WL_TK[23] WL_TK[24] WL_TK[25] WL_TK[26] WL_TK[27] WL_TK[28] WL_TK[29] 
+ WL_TK[30] WL_TK[31] NET60[0] NET60[1] NET60[2] NET60[3] NET60[4] NET60[5] 
+ NET60[6] NET60[7] NET59 NET69 NET57[0] NET57[1] NET57[2] NET57[3] NET57[4] 
+ NET57[5] NET57[6] NET57[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
XTRKNORX16_DUMY1 BL_TK VDDI VSSI WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] 
+ WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] 
+ WL_TK[32] WL_TK[33] WL_TK[34] WL_TK[35] WL_TK[36] WL_TK[37] WL_TK[38] 
+ WL_TK[39] WL_TK[40] WL_TK[41] WL_TK[42] WL_TK[43] WL_TK[44] WL_TK[45] 
+ WL_TK[46] WL_TK[47] NET50[0] NET50[1] NET50[2] NET50[3] NET50[4] NET50[5] 
+ NET50[6] NET50[7] NET49 NET59 NET47[0] NET47[1] NET47[2] NET47[3] NET47[4] 
+ NET47[5] NET47[6] NET47[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
XTRKNORX16_BCELL BL_TK VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] 
+ WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL_TK[0] 
+ WL_TK[1] WL_TK[2] WL_TK[3] WL_TK[4] WL_TK[5] WL_TK[6] WL_TK[7] WL_TK[8] 
+ WL_TK[9] WL_TK[10] WL_TK[11] WL_TK[12] WL_TK[13] WL_TK[14] WL_TK[15] 
+ NET70[0] NET70[1] NET70[2] NET70[3] NET70[4] NET70[5] NET70[6] NET70[7] 
+ NET69 NET68 NET67[0] NET67[1] NET67[2] NET67[3] NET67[4] NET67[5] NET67[6] 
+ NET67[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
XTRKNORX16_DUMY2 BL_TK VDDI VSSI WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] 
+ WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] 
+ WL_TK[48] WL_TK[49] WL_TK[50] WL_TK[51] WL_TK[52] WL_TK[53] WL_TK[54] 
+ WL_TK[55] WL_TK[56] WL_TK[57] WL_TK[58] WL_TK[59] WL_TK[60] WL_TK[61] 
+ WL_TK[62] WL_TK[63] NET40[0] NET40[1] NET40[2] NET40[3] NET40[4] NET40[5] 
+ NET40[6] NET40[7] NET39 NET49 NET37[0] NET37[1] NET37[2] NET37[3] NET37[4] 
+ NET37[5] NET37[6] NET37[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    TKBL_S16_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TKBL_S16_CHAR BL_TK VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL_TK[0] 
+ WL_TK[1] WL_TK[2] WL_TK[3] WL_TK[4] WL_TK[5] WL_TK[6] WL_TK[7] WL_TK[8] 
+ WL_TK[9] WL_TK[10] WL_TK[11] WL_TK[12] WL_TK[13] WL_TK[14] WL_TK[15] TIEH 
+ TIEL
*.PININFO BL_TK:B VDDI:B VSSI:B WL[0]:B WL[1]:B WL[2]:B WL[3]:B WL[4]:B 
*.PININFO WL[5]:B WL[6]:B WL[7]:B WL[8]:B WL[9]:B WL[10]:B WL[11]:B WL[12]:B 
*.PININFO WL[13]:B WL[14]:B WL[15]:B WL_TK[0]:B WL_TK[1]:B WL_TK[2]:B 
*.PININFO WL_TK[3]:B WL_TK[4]:B WL_TK[5]:B WL_TK[6]:B WL_TK[7]:B WL_TK[8]:B 
*.PININFO WL_TK[9]:B WL_TK[10]:B WL_TK[11]:B WL_TK[12]:B WL_TK[13]:B 
*.PININFO WL_TK[14]:B WL_TK[15]:B TIEH:B TIEL:B
XTRKNORX16_BCELL BL_TK VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] 
+ WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL_TK[0] 
+ WL_TK[1] WL_TK[2] WL_TK[3] WL_TK[4] WL_TK[5] WL_TK[6] WL_TK[7] WL_TK[8] 
+ WL_TK[9] WL_TK[10] WL_TK[11] WL_TK[12] WL_TK[13] WL_TK[14] WL_TK[15] 
+ NET70[0] NET70[1] NET70[2] NET70[3] NET70[4] NET70[5] NET70[6] NET70[7] 
+ NET69 NET68 NET67[0] NET67[1] NET67[2] NET67[3] NET67[4] NET67[5] NET67[6] 
+ NET67[7] TIEH S1AHSF400W40_TRKNORX16_CHAR
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    TKBL_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TKBL_SIM BL_TK_BT BL_TK_TP CVDDHD PD VDDHD VDDI VSSI WL[0] WL[1] WL[2] 
+ WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] 
+ WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] 
+ WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] 
+ WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] 
+ WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] 
+ WL[59] WL[60] WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] 
+ WL[70] WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] 
+ WL[81] WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] 
+ WL[92] WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] 
+ WL[102] WL[103] WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] 
+ WL[111] WL[112] WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] 
+ WL[120] WL[121] WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] 
+ WL[129] WL[130] WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] 
+ WL[138] WL[139] WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] 
+ WL[147] WL[148] WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] 
+ WL[156] WL[157] WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] 
+ WL[165] WL[166] WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] 
+ WL[174] WL[175] WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] 
+ WL[183] WL[184] WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] 
+ WL[192] WL[193] WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] 
+ WL[201] WL[202] WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] 
+ WL[210] WL[211] WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] 
+ WL[219] WL[220] WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] 
+ WL[228] WL[229] WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] 
+ WL[237] WL[238] WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] 
+ WL[246] WL[247] WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] 
+ WL[255] WL[256] WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] 
+ WL[264] WL[265] WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] 
+ WL[273] WL[274] WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] 
+ WL[282] WL[283] WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] 
+ WL[291] WL[292] WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] 
+ WL[300] WL[301] WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] 
+ WL[309] WL[310] WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] 
+ WL[318] WL[319] WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] 
+ WL[327] WL[328] WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] 
+ WL[336] WL[337] WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] 
+ WL[345] WL[346] WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] 
+ WL[354] WL[355] WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] 
+ WL[363] WL[364] WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] 
+ WL[372] WL[373] WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] 
+ WL[381] WL[382] WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] 
+ WL[390] WL[391] WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] 
+ WL[399] WL[400] WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] 
+ WL[408] WL[409] WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] 
+ WL[417] WL[418] WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] 
+ WL[426] WL[427] WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] 
+ WL[435] WL[436] WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] 
+ WL[444] WL[445] WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] 
+ WL[453] WL[454] WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] 
+ WL[462] WL[463] WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] 
+ WL[471] WL[472] WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] 
+ WL[480] WL[481] WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] 
+ WL[489] WL[490] WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] 
+ WL[498] WL[499] WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] 
+ WL[507] WL[508] WL[509] WL[510] WL[511] WL_TK[0] WL_TK[1] WL_TK[2] WL_TK[3] 
+ WL_TK[4] WL_TK[5] WL_TK[6] WL_TK[7] WL_TK[8] WL_TK[9] WL_TK[10] WL_TK[11] 
+ WL_TK[12] WL_TK[13] WL_TK[14] WL_TK[15] WL_TK[16] WL_TK[17] WL_TK[18] 
+ WL_TK[19] WL_TK[20] WL_TK[21] WL_TK[22] WL_TK[23] WL_TK[24] WL_TK[25] 
+ WL_TK[26] WL_TK[27] WL_TK[28] WL_TK[29] WL_TK[30] WL_TK[31] WL_TK[32] 
+ WL_TK[33] WL_TK[34] WL_TK[35] WL_TK[36] WL_TK[37] WL_TK[38] WL_TK[39] 
+ WL_TK[40] WL_TK[41] WL_TK[42] WL_TK[43] WL_TK[44] WL_TK[45] WL_TK[46] 
+ WL_TK[47] WL_TK[48] WL_TK[49] WL_TK[50] WL_TK[51] WL_TK[52] WL_TK[53] 
+ WL_TK[54] WL_TK[55] WL_TK[56] WL_TK[57] WL_TK[58] WL_TK[59] WL_TK[60] 
+ WL_TK[61] WL_TK[62] WL_TK[63] WL_TK[64] WL_TK[65] WL_TK[66] WL_TK[67] 
+ WL_TK[68] WL_TK[69] WL_TK[70] WL_TK[71] WL_TK[72] WL_TK[73] WL_TK[74] 
+ WL_TK[75] WL_TK[76] WL_TK[77] WL_TK[78] WL_TK[79] WL_TK[80] WL_TK[81] 
+ WL_TK[82] WL_TK[83] WL_TK[84] WL_TK[85] WL_TK[86] WL_TK[87] WL_TK[88] 
+ WL_TK[89] WL_TK[90] WL_TK[91] WL_TK[92] WL_TK[93] WL_TK[94] WL_TK[95] 
+ WL_TK[96] WL_TK[97] WL_TK[98] WL_TK[99] WL_TK[100] WL_TK[101] WL_TK[102] 
+ WL_TK[103] WL_TK[104] WL_TK[105] WL_TK[106] WL_TK[107] WL_TK[108] WL_TK[109] 
+ WL_TK[110] WL_TK[111] WL_TK[112] WL_TK[113] WL_TK[114] WL_TK[115] WL_TK[116] 
+ WL_TK[117] WL_TK[118] WL_TK[119] WL_TK[120] WL_TK[121] WL_TK[122] WL_TK[123] 
+ WL_TK[124] WL_TK[125] WL_TK[126] WL_TK[127] WL_TK[128] WL_TK[129] WL_TK[130] 
+ WL_TK[131] WL_TK[132] WL_TK[133] WL_TK[134] WL_TK[135] WL_TK[136] WL_TK[137] 
+ WL_TK[138] WL_TK[139] WL_TK[140] WL_TK[141] WL_TK[142] WL_TK[143] WL_TK[144] 
+ WL_TK[145] WL_TK[146] WL_TK[147] WL_TK[148] WL_TK[149] WL_TK[150] WL_TK[151] 
+ WL_TK[152] WL_TK[153] WL_TK[154] WL_TK[155] WL_TK[156] WL_TK[157] WL_TK[158] 
+ WL_TK[159] WL_TK[160] WL_TK[161] WL_TK[162] WL_TK[163] WL_TK[164] WL_TK[165] 
+ WL_TK[166] WL_TK[167] WL_TK[168] WL_TK[169] WL_TK[170] WL_TK[171] WL_TK[172] 
+ WL_TK[173] WL_TK[174] WL_TK[175] WL_TK[176] WL_TK[177] WL_TK[178] WL_TK[179] 
+ WL_TK[180] WL_TK[181] WL_TK[182] WL_TK[183] WL_TK[184] WL_TK[185] WL_TK[186] 
+ WL_TK[187] WL_TK[188] WL_TK[189] WL_TK[190] WL_TK[191] WL_TK[192] WL_TK[193] 
+ WL_TK[194] WL_TK[195] WL_TK[196] WL_TK[197] WL_TK[198] WL_TK[199] WL_TK[200] 
+ WL_TK[201] WL_TK[202] WL_TK[203] WL_TK[204] WL_TK[205] WL_TK[206] WL_TK[207] 
+ WL_TK[208] WL_TK[209] WL_TK[210] WL_TK[211] WL_TK[212] WL_TK[213] WL_TK[214] 
+ WL_TK[215] WL_TK[216] WL_TK[217] WL_TK[218] WL_TK[219] WL_TK[220] WL_TK[221] 
+ WL_TK[222] WL_TK[223] WL_TK[224] WL_TK[225] WL_TK[226] WL_TK[227] WL_TK[228] 
+ WL_TK[229] WL_TK[230] WL_TK[231] WL_TK[232] WL_TK[233] WL_TK[234] WL_TK[235] 
+ WL_TK[236] WL_TK[237] WL_TK[238] WL_TK[239] WL_TK[240] WL_TK[241] WL_TK[242] 
+ WL_TK[243] WL_TK[244] WL_TK[245] WL_TK[246] WL_TK[247] WL_TK[248] WL_TK[249] 
+ WL_TK[250] WL_TK[251] WL_TK[252] WL_TK[253] WL_TK[254] WL_TK[255] WL_TK[256] 
+ WL_TK[257] WL_TK[258] WL_TK[259] WL_TK[260] WL_TK[261] WL_TK[262] WL_TK[263] 
+ WL_TK[264] WL_TK[265] WL_TK[266] WL_TK[267] WL_TK[268] WL_TK[269] WL_TK[270] 
+ WL_TK[271] WL_TK[272] WL_TK[273] WL_TK[274] WL_TK[275] WL_TK[276] WL_TK[277] 
+ WL_TK[278] WL_TK[279] WL_TK[280] WL_TK[281] WL_TK[282] WL_TK[283] WL_TK[284] 
+ WL_TK[285] WL_TK[286] WL_TK[287] WL_TK[288] WL_TK[289] WL_TK[290] WL_TK[291] 
+ WL_TK[292] WL_TK[293] WL_TK[294] WL_TK[295] WL_TK[296] WL_TK[297] WL_TK[298] 
+ WL_TK[299] WL_TK[300] WL_TK[301] WL_TK[302] WL_TK[303] WL_TK[304] WL_TK[305] 
+ WL_TK[306] WL_TK[307] WL_TK[308] WL_TK[309] WL_TK[310] WL_TK[311] WL_TK[312] 
+ WL_TK[313] WL_TK[314] WL_TK[315] WL_TK[316] WL_TK[317] WL_TK[318] WL_TK[319] 
+ WL_TK[320] WL_TK[321] WL_TK[322] WL_TK[323] WL_TK[324] WL_TK[325] WL_TK[326] 
+ WL_TK[327] WL_TK[328] WL_TK[329] WL_TK[330] WL_TK[331] WL_TK[332] WL_TK[333] 
+ WL_TK[334] WL_TK[335] WL_TK[336] WL_TK[337] WL_TK[338] WL_TK[339] WL_TK[340] 
+ WL_TK[341] WL_TK[342] WL_TK[343] WL_TK[344] WL_TK[345] WL_TK[346] WL_TK[347] 
+ WL_TK[348] WL_TK[349] WL_TK[350] WL_TK[351] WL_TK[352] WL_TK[353] WL_TK[354] 
+ WL_TK[355] WL_TK[356] WL_TK[357] WL_TK[358] WL_TK[359] WL_TK[360] WL_TK[361] 
+ WL_TK[362] WL_TK[363] WL_TK[364] WL_TK[365] WL_TK[366] WL_TK[367] WL_TK[368] 
+ WL_TK[369] WL_TK[370] WL_TK[371] WL_TK[372] WL_TK[373] WL_TK[374] WL_TK[375] 
+ WL_TK[376] WL_TK[377] WL_TK[378] WL_TK[379] WL_TK[380] WL_TK[381] WL_TK[382] 
+ WL_TK[383] WL_TK[384] WL_TK[385] WL_TK[386] WL_TK[387] WL_TK[388] WL_TK[389] 
+ WL_TK[390] WL_TK[391] WL_TK[392] WL_TK[393] WL_TK[394] WL_TK[395] WL_TK[396] 
+ WL_TK[397] WL_TK[398] WL_TK[399] WL_TK[400] WL_TK[401] WL_TK[402] WL_TK[403] 
+ WL_TK[404] WL_TK[405] WL_TK[406] WL_TK[407] WL_TK[408] WL_TK[409] WL_TK[410] 
+ WL_TK[411] WL_TK[412] WL_TK[413] WL_TK[414] WL_TK[415] WL_TK[416] WL_TK[417] 
+ WL_TK[418] WL_TK[419] WL_TK[420] WL_TK[421] WL_TK[422] WL_TK[423] WL_TK[424] 
+ WL_TK[425] WL_TK[426] WL_TK[427] WL_TK[428] WL_TK[429] WL_TK[430] WL_TK[431] 
+ WL_TK[432] WL_TK[433] WL_TK[434] WL_TK[435] WL_TK[436] WL_TK[437] WL_TK[438] 
+ WL_TK[439] WL_TK[440] WL_TK[441] WL_TK[442] WL_TK[443] WL_TK[444] WL_TK[445] 
+ WL_TK[446] WL_TK[447] WL_TK[448] WL_TK[449] WL_TK[450] WL_TK[451] WL_TK[452] 
+ WL_TK[453] WL_TK[454] WL_TK[455] WL_TK[456] WL_TK[457] WL_TK[458] WL_TK[459] 
+ WL_TK[460] WL_TK[461] WL_TK[462] WL_TK[463] WL_TK[464] WL_TK[465] WL_TK[466] 
+ WL_TK[467] WL_TK[468] WL_TK[469] WL_TK[470] WL_TK[471] WL_TK[472] WL_TK[473] 
+ WL_TK[474] WL_TK[475] WL_TK[476] WL_TK[477] WL_TK[478] WL_TK[479] WL_TK[480] 
+ WL_TK[481] WL_TK[482] WL_TK[483] WL_TK[484] WL_TK[485] WL_TK[486] WL_TK[487] 
+ WL_TK[488] WL_TK[489] WL_TK[490] WL_TK[491] WL_TK[492] WL_TK[493] WL_TK[494] 
+ WL_TK[495] WL_TK[496] WL_TK[497] WL_TK[498] WL_TK[499] WL_TK[500] WL_TK[501] 
+ WL_TK[502] WL_TK[503] WL_TK[504] WL_TK[505] WL_TK[506] WL_TK[507] WL_TK[508] 
+ WL_TK[509] WL_TK[510] WL_TK[511] TIEH TIEL
*.PININFO PD:I BL_TK_BT:B BL_TK_TP:B CVDDHD:B VDDHD:B VDDI:B VSSI:B WL[0]:B 
*.PININFO WL[1]:B WL[2]:B WL[3]:B WL[4]:B WL[5]:B WL[6]:B WL[7]:B WL[8]:B 
*.PININFO WL[9]:B WL[10]:B WL[11]:B WL[12]:B WL[13]:B WL[14]:B WL[15]:B 
*.PININFO WL[16]:B WL[17]:B WL[18]:B WL[19]:B WL[20]:B WL[21]:B WL[22]:B 
*.PININFO WL[23]:B WL[24]:B WL[25]:B WL[26]:B WL[27]:B WL[28]:B WL[29]:B 
*.PININFO WL[30]:B WL[31]:B WL[32]:B WL[33]:B WL[34]:B WL[35]:B WL[36]:B 
*.PININFO WL[37]:B WL[38]:B WL[39]:B WL[40]:B WL[41]:B WL[42]:B WL[43]:B 
*.PININFO WL[44]:B WL[45]:B WL[46]:B WL[47]:B WL[48]:B WL[49]:B WL[50]:B 
*.PININFO WL[51]:B WL[52]:B WL[53]:B WL[54]:B WL[55]:B WL[56]:B WL[57]:B 
*.PININFO WL[58]:B WL[59]:B WL[60]:B WL[61]:B WL[62]:B WL[63]:B WL[64]:B 
*.PININFO WL[65]:B WL[66]:B WL[67]:B WL[68]:B WL[69]:B WL[70]:B WL[71]:B 
*.PININFO WL[72]:B WL[73]:B WL[74]:B WL[75]:B WL[76]:B WL[77]:B WL[78]:B 
*.PININFO WL[79]:B WL[80]:B WL[81]:B WL[82]:B WL[83]:B WL[84]:B WL[85]:B 
*.PININFO WL[86]:B WL[87]:B WL[88]:B WL[89]:B WL[90]:B WL[91]:B WL[92]:B 
*.PININFO WL[93]:B WL[94]:B WL[95]:B WL[96]:B WL[97]:B WL[98]:B WL[99]:B 
*.PININFO WL[100]:B WL[101]:B WL[102]:B WL[103]:B WL[104]:B WL[105]:B 
*.PININFO WL[106]:B WL[107]:B WL[108]:B WL[109]:B WL[110]:B WL[111]:B 
*.PININFO WL[112]:B WL[113]:B WL[114]:B WL[115]:B WL[116]:B WL[117]:B 
*.PININFO WL[118]:B WL[119]:B WL[120]:B WL[121]:B WL[122]:B WL[123]:B 
*.PININFO WL[124]:B WL[125]:B WL[126]:B WL[127]:B WL[128]:B WL[129]:B 
*.PININFO WL[130]:B WL[131]:B WL[132]:B WL[133]:B WL[134]:B WL[135]:B 
*.PININFO WL[136]:B WL[137]:B WL[138]:B WL[139]:B WL[140]:B WL[141]:B 
*.PININFO WL[142]:B WL[143]:B WL[144]:B WL[145]:B WL[146]:B WL[147]:B 
*.PININFO WL[148]:B WL[149]:B WL[150]:B WL[151]:B WL[152]:B WL[153]:B 
*.PININFO WL[154]:B WL[155]:B WL[156]:B WL[157]:B WL[158]:B WL[159]:B 
*.PININFO WL[160]:B WL[161]:B WL[162]:B WL[163]:B WL[164]:B WL[165]:B 
*.PININFO WL[166]:B WL[167]:B WL[168]:B WL[169]:B WL[170]:B WL[171]:B 
*.PININFO WL[172]:B WL[173]:B WL[174]:B WL[175]:B WL[176]:B WL[177]:B 
*.PININFO WL[178]:B WL[179]:B WL[180]:B WL[181]:B WL[182]:B WL[183]:B 
*.PININFO WL[184]:B WL[185]:B WL[186]:B WL[187]:B WL[188]:B WL[189]:B 
*.PININFO WL[190]:B WL[191]:B WL[192]:B WL[193]:B WL[194]:B WL[195]:B 
*.PININFO WL[196]:B WL[197]:B WL[198]:B WL[199]:B WL[200]:B WL[201]:B 
*.PININFO WL[202]:B WL[203]:B WL[204]:B WL[205]:B WL[206]:B WL[207]:B 
*.PININFO WL[208]:B WL[209]:B WL[210]:B WL[211]:B WL[212]:B WL[213]:B 
*.PININFO WL[214]:B WL[215]:B WL[216]:B WL[217]:B WL[218]:B WL[219]:B 
*.PININFO WL[220]:B WL[221]:B WL[222]:B WL[223]:B WL[224]:B WL[225]:B 
*.PININFO WL[226]:B WL[227]:B WL[228]:B WL[229]:B WL[230]:B WL[231]:B 
*.PININFO WL[232]:B WL[233]:B WL[234]:B WL[235]:B WL[236]:B WL[237]:B 
*.PININFO WL[238]:B WL[239]:B WL[240]:B WL[241]:B WL[242]:B WL[243]:B 
*.PININFO WL[244]:B WL[245]:B WL[246]:B WL[247]:B WL[248]:B WL[249]:B 
*.PININFO WL[250]:B WL[251]:B WL[252]:B WL[253]:B WL[254]:B WL[255]:B 
*.PININFO WL[256]:B WL[257]:B WL[258]:B WL[259]:B WL[260]:B WL[261]:B 
*.PININFO WL[262]:B WL[263]:B WL[264]:B WL[265]:B WL[266]:B WL[267]:B 
*.PININFO WL[268]:B WL[269]:B WL[270]:B WL[271]:B WL[272]:B WL[273]:B 
*.PININFO WL[274]:B WL[275]:B WL[276]:B WL[277]:B WL[278]:B WL[279]:B 
*.PININFO WL[280]:B WL[281]:B WL[282]:B WL[283]:B WL[284]:B WL[285]:B 
*.PININFO WL[286]:B WL[287]:B WL[288]:B WL[289]:B WL[290]:B WL[291]:B 
*.PININFO WL[292]:B WL[293]:B WL[294]:B WL[295]:B WL[296]:B WL[297]:B 
*.PININFO WL[298]:B WL[299]:B WL[300]:B WL[301]:B WL[302]:B WL[303]:B 
*.PININFO WL[304]:B WL[305]:B WL[306]:B WL[307]:B WL[308]:B WL[309]:B 
*.PININFO WL[310]:B WL[311]:B WL[312]:B WL[313]:B WL[314]:B WL[315]:B 
*.PININFO WL[316]:B WL[317]:B WL[318]:B WL[319]:B WL[320]:B WL[321]:B 
*.PININFO WL[322]:B WL[323]:B WL[324]:B WL[325]:B WL[326]:B WL[327]:B 
*.PININFO WL[328]:B WL[329]:B WL[330]:B WL[331]:B WL[332]:B WL[333]:B 
*.PININFO WL[334]:B WL[335]:B WL[336]:B WL[337]:B WL[338]:B WL[339]:B 
*.PININFO WL[340]:B WL[341]:B WL[342]:B WL[343]:B WL[344]:B WL[345]:B 
*.PININFO WL[346]:B WL[347]:B WL[348]:B WL[349]:B WL[350]:B WL[351]:B 
*.PININFO WL[352]:B WL[353]:B WL[354]:B WL[355]:B WL[356]:B WL[357]:B 
*.PININFO WL[358]:B WL[359]:B WL[360]:B WL[361]:B WL[362]:B WL[363]:B 
*.PININFO WL[364]:B WL[365]:B WL[366]:B WL[367]:B WL[368]:B WL[369]:B 
*.PININFO WL[370]:B WL[371]:B WL[372]:B WL[373]:B WL[374]:B WL[375]:B 
*.PININFO WL[376]:B WL[377]:B WL[378]:B WL[379]:B WL[380]:B WL[381]:B 
*.PININFO WL[382]:B WL[383]:B WL[384]:B WL[385]:B WL[386]:B WL[387]:B 
*.PININFO WL[388]:B WL[389]:B WL[390]:B WL[391]:B WL[392]:B WL[393]:B 
*.PININFO WL[394]:B WL[395]:B WL[396]:B WL[397]:B WL[398]:B WL[399]:B 
*.PININFO WL[400]:B WL[401]:B WL[402]:B WL[403]:B WL[404]:B WL[405]:B 
*.PININFO WL[406]:B WL[407]:B WL[408]:B WL[409]:B WL[410]:B WL[411]:B 
*.PININFO WL[412]:B WL[413]:B WL[414]:B WL[415]:B WL[416]:B WL[417]:B 
*.PININFO WL[418]:B WL[419]:B WL[420]:B WL[421]:B WL[422]:B WL[423]:B 
*.PININFO WL[424]:B WL[425]:B WL[426]:B WL[427]:B WL[428]:B WL[429]:B 
*.PININFO WL[430]:B WL[431]:B WL[432]:B WL[433]:B WL[434]:B WL[435]:B 
*.PININFO WL[436]:B WL[437]:B WL[438]:B WL[439]:B WL[440]:B WL[441]:B 
*.PININFO WL[442]:B WL[443]:B WL[444]:B WL[445]:B WL[446]:B WL[447]:B 
*.PININFO WL[448]:B WL[449]:B WL[450]:B WL[451]:B WL[452]:B WL[453]:B 
*.PININFO WL[454]:B WL[455]:B WL[456]:B WL[457]:B WL[458]:B WL[459]:B 
*.PININFO WL[460]:B WL[461]:B WL[462]:B WL[463]:B WL[464]:B WL[465]:B 
*.PININFO WL[466]:B WL[467]:B WL[468]:B WL[469]:B WL[470]:B WL[471]:B 
*.PININFO WL[472]:B WL[473]:B WL[474]:B WL[475]:B WL[476]:B WL[477]:B 
*.PININFO WL[478]:B WL[479]:B WL[480]:B WL[481]:B WL[482]:B WL[483]:B 
*.PININFO WL[484]:B WL[485]:B WL[486]:B WL[487]:B WL[488]:B WL[489]:B 
*.PININFO WL[490]:B WL[491]:B WL[492]:B WL[493]:B WL[494]:B WL[495]:B 
*.PININFO WL[496]:B WL[497]:B WL[498]:B WL[499]:B WL[500]:B WL[501]:B 
*.PININFO WL[502]:B WL[503]:B WL[504]:B WL[505]:B WL[506]:B WL[507]:B 
*.PININFO WL[508]:B WL[509]:B WL[510]:B WL[511]:B WL_TK[0]:B WL_TK[1]:B 
*.PININFO WL_TK[2]:B WL_TK[3]:B WL_TK[4]:B WL_TK[5]:B WL_TK[6]:B WL_TK[7]:B 
*.PININFO WL_TK[8]:B WL_TK[9]:B WL_TK[10]:B WL_TK[11]:B WL_TK[12]:B 
*.PININFO WL_TK[13]:B WL_TK[14]:B WL_TK[15]:B WL_TK[16]:B WL_TK[17]:B 
*.PININFO WL_TK[18]:B WL_TK[19]:B WL_TK[20]:B WL_TK[21]:B WL_TK[22]:B 
*.PININFO WL_TK[23]:B WL_TK[24]:B WL_TK[25]:B WL_TK[26]:B WL_TK[27]:B 
*.PININFO WL_TK[28]:B WL_TK[29]:B WL_TK[30]:B WL_TK[31]:B WL_TK[32]:B 
*.PININFO WL_TK[33]:B WL_TK[34]:B WL_TK[35]:B WL_TK[36]:B WL_TK[37]:B 
*.PININFO WL_TK[38]:B WL_TK[39]:B WL_TK[40]:B WL_TK[41]:B WL_TK[42]:B 
*.PININFO WL_TK[43]:B WL_TK[44]:B WL_TK[45]:B WL_TK[46]:B WL_TK[47]:B 
*.PININFO WL_TK[48]:B WL_TK[49]:B WL_TK[50]:B WL_TK[51]:B WL_TK[52]:B 
*.PININFO WL_TK[53]:B WL_TK[54]:B WL_TK[55]:B WL_TK[56]:B WL_TK[57]:B 
*.PININFO WL_TK[58]:B WL_TK[59]:B WL_TK[60]:B WL_TK[61]:B WL_TK[62]:B 
*.PININFO WL_TK[63]:B WL_TK[64]:B WL_TK[65]:B WL_TK[66]:B WL_TK[67]:B 
*.PININFO WL_TK[68]:B WL_TK[69]:B WL_TK[70]:B WL_TK[71]:B WL_TK[72]:B 
*.PININFO WL_TK[73]:B WL_TK[74]:B WL_TK[75]:B WL_TK[76]:B WL_TK[77]:B 
*.PININFO WL_TK[78]:B WL_TK[79]:B WL_TK[80]:B WL_TK[81]:B WL_TK[82]:B 
*.PININFO WL_TK[83]:B WL_TK[84]:B WL_TK[85]:B WL_TK[86]:B WL_TK[87]:B 
*.PININFO WL_TK[88]:B WL_TK[89]:B WL_TK[90]:B WL_TK[91]:B WL_TK[92]:B 
*.PININFO WL_TK[93]:B WL_TK[94]:B WL_TK[95]:B WL_TK[96]:B WL_TK[97]:B 
*.PININFO WL_TK[98]:B WL_TK[99]:B WL_TK[100]:B WL_TK[101]:B WL_TK[102]:B 
*.PININFO WL_TK[103]:B WL_TK[104]:B WL_TK[105]:B WL_TK[106]:B WL_TK[107]:B 
*.PININFO WL_TK[108]:B WL_TK[109]:B WL_TK[110]:B WL_TK[111]:B WL_TK[112]:B 
*.PININFO WL_TK[113]:B WL_TK[114]:B WL_TK[115]:B WL_TK[116]:B WL_TK[117]:B 
*.PININFO WL_TK[118]:B WL_TK[119]:B WL_TK[120]:B WL_TK[121]:B WL_TK[122]:B 
*.PININFO WL_TK[123]:B WL_TK[124]:B WL_TK[125]:B WL_TK[126]:B WL_TK[127]:B 
*.PININFO WL_TK[128]:B WL_TK[129]:B WL_TK[130]:B WL_TK[131]:B WL_TK[132]:B 
*.PININFO WL_TK[133]:B WL_TK[134]:B WL_TK[135]:B WL_TK[136]:B WL_TK[137]:B 
*.PININFO WL_TK[138]:B WL_TK[139]:B WL_TK[140]:B WL_TK[141]:B WL_TK[142]:B 
*.PININFO WL_TK[143]:B WL_TK[144]:B WL_TK[145]:B WL_TK[146]:B WL_TK[147]:B 
*.PININFO WL_TK[148]:B WL_TK[149]:B WL_TK[150]:B WL_TK[151]:B WL_TK[152]:B 
*.PININFO WL_TK[153]:B WL_TK[154]:B WL_TK[155]:B WL_TK[156]:B WL_TK[157]:B 
*.PININFO WL_TK[158]:B WL_TK[159]:B WL_TK[160]:B WL_TK[161]:B WL_TK[162]:B 
*.PININFO WL_TK[163]:B WL_TK[164]:B WL_TK[165]:B WL_TK[166]:B WL_TK[167]:B 
*.PININFO WL_TK[168]:B WL_TK[169]:B WL_TK[170]:B WL_TK[171]:B WL_TK[172]:B 
*.PININFO WL_TK[173]:B WL_TK[174]:B WL_TK[175]:B WL_TK[176]:B WL_TK[177]:B 
*.PININFO WL_TK[178]:B WL_TK[179]:B WL_TK[180]:B WL_TK[181]:B WL_TK[182]:B 
*.PININFO WL_TK[183]:B WL_TK[184]:B WL_TK[185]:B WL_TK[186]:B WL_TK[187]:B 
*.PININFO WL_TK[188]:B WL_TK[189]:B WL_TK[190]:B WL_TK[191]:B WL_TK[192]:B 
*.PININFO WL_TK[193]:B WL_TK[194]:B WL_TK[195]:B WL_TK[196]:B WL_TK[197]:B 
*.PININFO WL_TK[198]:B WL_TK[199]:B WL_TK[200]:B WL_TK[201]:B WL_TK[202]:B 
*.PININFO WL_TK[203]:B WL_TK[204]:B WL_TK[205]:B WL_TK[206]:B WL_TK[207]:B 
*.PININFO WL_TK[208]:B WL_TK[209]:B WL_TK[210]:B WL_TK[211]:B WL_TK[212]:B 
*.PININFO WL_TK[213]:B WL_TK[214]:B WL_TK[215]:B WL_TK[216]:B WL_TK[217]:B 
*.PININFO WL_TK[218]:B WL_TK[219]:B WL_TK[220]:B WL_TK[221]:B WL_TK[222]:B 
*.PININFO WL_TK[223]:B WL_TK[224]:B WL_TK[225]:B WL_TK[226]:B WL_TK[227]:B 
*.PININFO WL_TK[228]:B WL_TK[229]:B WL_TK[230]:B WL_TK[231]:B WL_TK[232]:B 
*.PININFO WL_TK[233]:B WL_TK[234]:B WL_TK[235]:B WL_TK[236]:B WL_TK[237]:B 
*.PININFO WL_TK[238]:B WL_TK[239]:B WL_TK[240]:B WL_TK[241]:B WL_TK[242]:B 
*.PININFO WL_TK[243]:B WL_TK[244]:B WL_TK[245]:B WL_TK[246]:B WL_TK[247]:B 
*.PININFO WL_TK[248]:B WL_TK[249]:B WL_TK[250]:B WL_TK[251]:B WL_TK[252]:B 
*.PININFO WL_TK[253]:B WL_TK[254]:B WL_TK[255]:B WL_TK[256]:B WL_TK[257]:B 
*.PININFO WL_TK[258]:B WL_TK[259]:B WL_TK[260]:B WL_TK[261]:B WL_TK[262]:B 
*.PININFO WL_TK[263]:B WL_TK[264]:B WL_TK[265]:B WL_TK[266]:B WL_TK[267]:B 
*.PININFO WL_TK[268]:B WL_TK[269]:B WL_TK[270]:B WL_TK[271]:B WL_TK[272]:B 
*.PININFO WL_TK[273]:B WL_TK[274]:B WL_TK[275]:B WL_TK[276]:B WL_TK[277]:B 
*.PININFO WL_TK[278]:B WL_TK[279]:B WL_TK[280]:B WL_TK[281]:B WL_TK[282]:B 
*.PININFO WL_TK[283]:B WL_TK[284]:B WL_TK[285]:B WL_TK[286]:B WL_TK[287]:B 
*.PININFO WL_TK[288]:B WL_TK[289]:B WL_TK[290]:B WL_TK[291]:B WL_TK[292]:B 
*.PININFO WL_TK[293]:B WL_TK[294]:B WL_TK[295]:B WL_TK[296]:B WL_TK[297]:B 
*.PININFO WL_TK[298]:B WL_TK[299]:B WL_TK[300]:B WL_TK[301]:B WL_TK[302]:B 
*.PININFO WL_TK[303]:B WL_TK[304]:B WL_TK[305]:B WL_TK[306]:B WL_TK[307]:B 
*.PININFO WL_TK[308]:B WL_TK[309]:B WL_TK[310]:B WL_TK[311]:B WL_TK[312]:B 
*.PININFO WL_TK[313]:B WL_TK[314]:B WL_TK[315]:B WL_TK[316]:B WL_TK[317]:B 
*.PININFO WL_TK[318]:B WL_TK[319]:B WL_TK[320]:B WL_TK[321]:B WL_TK[322]:B 
*.PININFO WL_TK[323]:B WL_TK[324]:B WL_TK[325]:B WL_TK[326]:B WL_TK[327]:B 
*.PININFO WL_TK[328]:B WL_TK[329]:B WL_TK[330]:B WL_TK[331]:B WL_TK[332]:B 
*.PININFO WL_TK[333]:B WL_TK[334]:B WL_TK[335]:B WL_TK[336]:B WL_TK[337]:B 
*.PININFO WL_TK[338]:B WL_TK[339]:B WL_TK[340]:B WL_TK[341]:B WL_TK[342]:B 
*.PININFO WL_TK[343]:B WL_TK[344]:B WL_TK[345]:B WL_TK[346]:B WL_TK[347]:B 
*.PININFO WL_TK[348]:B WL_TK[349]:B WL_TK[350]:B WL_TK[351]:B WL_TK[352]:B 
*.PININFO WL_TK[353]:B WL_TK[354]:B WL_TK[355]:B WL_TK[356]:B WL_TK[357]:B 
*.PININFO WL_TK[358]:B WL_TK[359]:B WL_TK[360]:B WL_TK[361]:B WL_TK[362]:B 
*.PININFO WL_TK[363]:B WL_TK[364]:B WL_TK[365]:B WL_TK[366]:B WL_TK[367]:B 
*.PININFO WL_TK[368]:B WL_TK[369]:B WL_TK[370]:B WL_TK[371]:B WL_TK[372]:B 
*.PININFO WL_TK[373]:B WL_TK[374]:B WL_TK[375]:B WL_TK[376]:B WL_TK[377]:B 
*.PININFO WL_TK[378]:B WL_TK[379]:B WL_TK[380]:B WL_TK[381]:B WL_TK[382]:B 
*.PININFO WL_TK[383]:B WL_TK[384]:B WL_TK[385]:B WL_TK[386]:B WL_TK[387]:B 
*.PININFO WL_TK[388]:B WL_TK[389]:B WL_TK[390]:B WL_TK[391]:B WL_TK[392]:B 
*.PININFO WL_TK[393]:B WL_TK[394]:B WL_TK[395]:B WL_TK[396]:B WL_TK[397]:B 
*.PININFO WL_TK[398]:B WL_TK[399]:B WL_TK[400]:B WL_TK[401]:B WL_TK[402]:B 
*.PININFO WL_TK[403]:B WL_TK[404]:B WL_TK[405]:B WL_TK[406]:B WL_TK[407]:B 
*.PININFO WL_TK[408]:B WL_TK[409]:B WL_TK[410]:B WL_TK[411]:B WL_TK[412]:B 
*.PININFO WL_TK[413]:B WL_TK[414]:B WL_TK[415]:B WL_TK[416]:B WL_TK[417]:B 
*.PININFO WL_TK[418]:B WL_TK[419]:B WL_TK[420]:B WL_TK[421]:B WL_TK[422]:B 
*.PININFO WL_TK[423]:B WL_TK[424]:B WL_TK[425]:B WL_TK[426]:B WL_TK[427]:B 
*.PININFO WL_TK[428]:B WL_TK[429]:B WL_TK[430]:B WL_TK[431]:B WL_TK[432]:B 
*.PININFO WL_TK[433]:B WL_TK[434]:B WL_TK[435]:B WL_TK[436]:B WL_TK[437]:B 
*.PININFO WL_TK[438]:B WL_TK[439]:B WL_TK[440]:B WL_TK[441]:B WL_TK[442]:B 
*.PININFO WL_TK[443]:B WL_TK[444]:B WL_TK[445]:B WL_TK[446]:B WL_TK[447]:B 
*.PININFO WL_TK[448]:B WL_TK[449]:B WL_TK[450]:B WL_TK[451]:B WL_TK[452]:B 
*.PININFO WL_TK[453]:B WL_TK[454]:B WL_TK[455]:B WL_TK[456]:B WL_TK[457]:B 
*.PININFO WL_TK[458]:B WL_TK[459]:B WL_TK[460]:B WL_TK[461]:B WL_TK[462]:B 
*.PININFO WL_TK[463]:B WL_TK[464]:B WL_TK[465]:B WL_TK[466]:B WL_TK[467]:B 
*.PININFO WL_TK[468]:B WL_TK[469]:B WL_TK[470]:B WL_TK[471]:B WL_TK[472]:B 
*.PININFO WL_TK[473]:B WL_TK[474]:B WL_TK[475]:B WL_TK[476]:B WL_TK[477]:B 
*.PININFO WL_TK[478]:B WL_TK[479]:B WL_TK[480]:B WL_TK[481]:B WL_TK[482]:B 
*.PININFO WL_TK[483]:B WL_TK[484]:B WL_TK[485]:B WL_TK[486]:B WL_TK[487]:B 
*.PININFO WL_TK[488]:B WL_TK[489]:B WL_TK[490]:B WL_TK[491]:B WL_TK[492]:B 
*.PININFO WL_TK[493]:B WL_TK[494]:B WL_TK[495]:B WL_TK[496]:B WL_TK[497]:B 
*.PININFO WL_TK[498]:B WL_TK[499]:B WL_TK[500]:B WL_TK[501]:B WL_TK[502]:B 
*.PININFO WL_TK[503]:B WL_TK[504]:B WL_TK[505]:B WL_TK[506]:B WL_TK[507]:B 
*.PININFO WL_TK[508]:B WL_TK[509]:B WL_TK[510]:B WL_TK[511]:B TIEH:B TIEL:B
XI13 NET034 NET06 NET028 NET027[0] NET027[1] NET027[2] NET027[3] NET027[4] 
+ NET027[5] NET027[6] NET027[7] NET027[8] NET027[9] NET027[10] NET027[11] 
+ NET027[12] NET027[13] NET027[14] NET027[15] NET027[16] NET027[17] NET027[18] 
+ NET027[19] NET027[20] NET027[21] NET027[22] NET027[23] NET027[24] NET027[25] 
+ NET027[26] NET027[27] NET027[28] NET027[29] NET027[30] NET027[31] NET027[32] 
+ NET027[33] NET027[34] NET027[35] NET027[36] NET027[37] NET027[38] NET027[39] 
+ NET027[40] NET027[41] NET027[42] NET027[43] NET027[44] NET027[45] NET027[46] 
+ NET027[47] NET027[48] NET027[49] NET027[50] NET027[51] NET027[52] NET027[53] 
+ NET027[54] NET027[55] NET027[56] NET027[57] NET027[58] NET027[59] NET027[60] 
+ NET027[61] NET027[62] NET027[63] NET027[64] NET027[65] NET027[66] NET027[67] 
+ NET027[68] NET027[69] NET027[70] NET027[71] NET027[72] NET027[73] NET027[74] 
+ NET027[75] NET027[76] NET027[77] NET027[78] NET027[79] NET027[80] NET027[81] 
+ NET027[82] NET027[83] NET027[84] NET027[85] NET027[86] NET027[87] NET027[88] 
+ NET027[89] NET027[90] NET027[91] NET027[92] NET027[93] NET027[94] NET027[95] 
+ NET027[96] NET027[97] NET027[98] NET027[99] NET027[100] NET027[101] 
+ NET027[102] NET027[103] NET027[104] NET027[105] NET027[106] NET027[107] 
+ NET027[108] NET027[109] NET027[110] NET027[111] NET027[112] NET027[113] 
+ NET027[114] NET027[115] NET027[116] NET027[117] NET027[118] NET027[119] 
+ NET027[120] NET027[121] NET027[122] NET027[123] NET027[124] NET027[125] 
+ NET027[126] NET027[127] NET027[128] NET027[129] NET027[130] NET027[131] 
+ NET027[132] NET027[133] NET027[134] NET027[135] NET027[136] NET027[137] 
+ NET027[138] NET027[139] NET027[140] NET027[141] NET027[142] NET027[143] 
+ NET027[144] NET027[145] NET027[146] NET027[147] NET027[148] NET027[149] 
+ NET027[150] NET027[151] NET027[152] NET027[153] NET027[154] NET027[155] 
+ NET027[156] NET027[157] NET027[158] NET027[159] NET027[160] NET027[161] 
+ NET027[162] NET027[163] NET027[164] NET027[165] NET027[166] NET027[167] 
+ NET027[168] NET027[169] NET027[170] NET027[171] NET027[172] NET027[173] 
+ NET027[174] NET027[175] NET027[176] NET027[177] NET027[178] NET027[179] 
+ NET027[180] NET027[181] NET027[182] NET027[183] NET027[184] NET027[185] 
+ NET027[186] NET027[187] NET027[188] NET027[189] NET027[190] NET027[191] 
+ NET027[192] NET027[193] NET027[194] NET027[195] NET027[196] NET027[197] 
+ NET027[198] NET027[199] NET027[200] NET027[201] NET027[202] NET027[203] 
+ NET027[204] NET027[205] NET027[206] NET027[207] NET027[208] NET027[209] 
+ NET027[210] NET027[211] NET027[212] NET027[213] NET027[214] NET027[215] 
+ NET027[216] NET027[217] NET027[218] NET027[219] NET027[220] NET027[221] 
+ NET027[222] NET027[223] NET027[224] NET027[225] NET027[226] NET027[227] 
+ NET027[228] NET027[229] NET027[230] NET027[231] NET027[232] NET027[233] 
+ NET027[234] NET027[235] NET027[236] NET027[237] NET027[238] NET027[239] 
+ NET027[240] NET027[241] NET027[242] NET027[243] NET027[244] NET027[245] 
+ NET027[246] NET027[247] NET027[248] NET027[249] NET027[250] NET027[251] 
+ NET027[252] NET027[253] NET027[254] NET027[255] NET027[256] NET027[257] 
+ NET027[258] NET027[259] NET027[260] NET027[261] NET027[262] NET027[263] 
+ NET027[264] NET027[265] NET027[266] NET027[267] NET027[268] NET027[269] 
+ NET027[270] NET027[271] NET027[272] NET027[273] NET027[274] NET027[275] 
+ NET027[276] NET027[277] NET027[278] NET027[279] NET027[280] NET027[281] 
+ NET027[282] NET027[283] NET027[284] NET027[285] NET027[286] NET027[287] 
+ NET027[288] NET027[289] NET027[290] NET027[291] NET027[292] NET027[293] 
+ NET027[294] NET027[295] NET027[296] NET027[297] NET027[298] NET027[299] 
+ NET027[300] NET027[301] NET027[302] NET027[303] NET027[304] NET027[305] 
+ NET027[306] NET027[307] NET027[308] NET027[309] NET027[310] NET027[311] 
+ NET027[312] NET027[313] NET027[314] NET027[315] NET027[316] NET027[317] 
+ NET027[318] NET027[319] NET027[320] NET027[321] NET027[322] NET027[323] 
+ NET027[324] NET027[325] NET027[326] NET027[327] NET027[328] NET027[329] 
+ NET027[330] NET027[331] NET027[332] NET027[333] NET027[334] NET027[335] 
+ NET027[336] NET027[337] NET027[338] NET027[339] NET027[340] NET027[341] 
+ NET027[342] NET027[343] NET027[344] NET027[345] NET027[346] NET027[347] 
+ NET027[348] NET027[349] NET027[350] NET027[351] NET027[352] NET027[353] 
+ NET027[354] NET027[355] NET027[356] NET027[357] NET027[358] NET027[359] 
+ NET027[360] NET027[361] NET027[362] NET027[363] NET027[364] NET027[365] 
+ NET027[366] NET027[367] NET027[368] NET027[369] NET027[370] NET027[371] 
+ NET027[372] NET027[373] NET027[374] NET027[375] NET027[376] NET027[377] 
+ NET027[378] NET027[379] NET027[380] NET027[381] NET027[382] NET027[383] 
+ NET027[384] NET027[385] NET027[386] NET027[387] NET027[388] NET027[389] 
+ NET027[390] NET027[391] NET027[392] NET027[393] NET027[394] NET027[395] 
+ NET027[396] NET027[397] NET027[398] NET027[399] NET027[400] NET027[401] 
+ NET027[402] NET027[403] NET027[404] NET027[405] NET027[406] NET027[407] 
+ NET027[408] NET027[409] NET027[410] NET027[411] NET027[412] NET027[413] 
+ NET027[414] NET027[415] NET027[416] NET027[417] NET027[418] NET027[419] 
+ NET027[420] NET027[421] NET027[422] NET027[423] NET027[424] NET027[425] 
+ NET027[426] NET027[427] NET027[428] NET027[429] NET027[430] NET027[431] 
+ NET027[432] NET027[433] NET027[434] NET027[435] NET027[436] NET027[437] 
+ NET027[438] NET027[439] NET027[440] NET027[441] NET027[442] NET027[443] 
+ NET027[444] NET027[445] NET027[446] NET027[447] NET027[448] NET027[449] 
+ NET027[450] NET027[451] NET027[452] NET027[453] NET027[454] NET027[455] 
+ NET027[456] NET027[457] NET027[458] NET027[459] NET027[460] NET027[461] 
+ NET027[462] NET027[463] NET027[464] NET027[465] NET027[466] NET027[467] 
+ NET027[468] NET027[469] NET027[470] NET027[471] NET027[472] NET027[473] 
+ NET027[474] NET027[475] NET027[476] NET027[477] NET027[478] NET027[479] 
+ NET027[480] NET027[481] NET027[482] NET027[483] NET027[484] NET027[485] 
+ NET027[486] NET027[487] NET027[488] NET027[489] NET027[490] NET027[491] 
+ NET027[492] NET027[493] NET027[494] NET027[495] NET027[496] NET027[497] 
+ NET027[498] NET027[499] NET027[500] NET027[501] NET027[502] NET027[503] 
+ NET027[504] NET027[505] NET027[506] NET027[507] NET027[508] NET027[509] 
+ NET027[510] NET027[511] NET05[0] NET05[1] NET05[2] NET05[3] NET05[4] 
+ NET05[5] NET05[6] NET05[7] NET05[8] NET05[9] NET05[10] NET05[11] NET05[12] 
+ NET05[13] NET05[14] NET05[15] NET05[16] NET05[17] NET05[18] NET05[19] 
+ NET05[20] NET05[21] NET05[22] NET05[23] NET05[24] NET05[25] NET05[26] 
+ NET05[27] NET05[28] NET05[29] NET05[30] NET05[31] NET05[32] NET05[33] 
+ NET05[34] NET05[35] NET05[36] NET05[37] NET05[38] NET05[39] NET05[40] 
+ NET05[41] NET05[42] NET05[43] NET05[44] NET05[45] NET05[46] NET05[47] 
+ NET05[48] NET05[49] NET05[50] NET05[51] NET05[52] NET05[53] NET05[54] 
+ NET05[55] NET05[56] NET05[57] NET05[58] NET05[59] NET05[60] NET05[61] 
+ NET05[62] NET05[63] NET05[64] NET05[65] NET05[66] NET05[67] NET05[68] 
+ NET05[69] NET05[70] NET05[71] NET05[72] NET05[73] NET05[74] NET05[75] 
+ NET05[76] NET05[77] NET05[78] NET05[79] NET05[80] NET05[81] NET05[82] 
+ NET05[83] NET05[84] NET05[85] NET05[86] NET05[87] NET05[88] NET05[89] 
+ NET05[90] NET05[91] NET05[92] NET05[93] NET05[94] NET05[95] NET05[96] 
+ NET05[97] NET05[98] NET05[99] NET05[100] NET05[101] NET05[102] NET05[103] 
+ NET05[104] NET05[105] NET05[106] NET05[107] NET05[108] NET05[109] NET05[110] 
+ NET05[111] NET05[112] NET05[113] NET05[114] NET05[115] NET05[116] NET05[117] 
+ NET05[118] NET05[119] NET05[120] NET05[121] NET05[122] NET05[123] NET05[124] 
+ NET05[125] NET05[126] NET05[127] NET05[128] NET05[129] NET05[130] NET05[131] 
+ NET05[132] NET05[133] NET05[134] NET05[135] NET05[136] NET05[137] NET05[138] 
+ NET05[139] NET05[140] NET05[141] NET05[142] NET05[143] NET05[144] NET05[145] 
+ NET05[146] NET05[147] NET05[148] NET05[149] NET05[150] NET05[151] NET05[152] 
+ NET05[153] NET05[154] NET05[155] NET05[156] NET05[157] NET05[158] NET05[159] 
+ NET05[160] NET05[161] NET05[162] NET05[163] NET05[164] NET05[165] NET05[166] 
+ NET05[167] NET05[168] NET05[169] NET05[170] NET05[171] NET05[172] NET05[173] 
+ NET05[174] NET05[175] NET05[176] NET05[177] NET05[178] NET05[179] NET05[180] 
+ NET05[181] NET05[182] NET05[183] NET05[184] NET05[185] NET05[186] NET05[187] 
+ NET05[188] NET05[189] NET05[190] NET05[191] NET05[192] NET05[193] NET05[194] 
+ NET05[195] NET05[196] NET05[197] NET05[198] NET05[199] NET05[200] NET05[201] 
+ NET05[202] NET05[203] NET05[204] NET05[205] NET05[206] NET05[207] NET05[208] 
+ NET05[209] NET05[210] NET05[211] NET05[212] NET05[213] NET05[214] NET05[215] 
+ NET05[216] NET05[217] NET05[218] NET05[219] NET05[220] NET05[221] NET05[222] 
+ NET05[223] NET05[224] NET05[225] NET05[226] NET05[227] NET05[228] NET05[229] 
+ NET05[230] NET05[231] NET05[232] NET05[233] NET05[234] NET05[235] NET05[236] 
+ NET05[237] NET05[238] NET05[239] NET05[240] NET05[241] NET05[242] NET05[243] 
+ NET05[244] NET05[245] NET05[246] NET05[247] NET05[248] NET05[249] NET05[250] 
+ NET05[251] NET05[252] NET05[253] NET05[254] NET05[255] NET05[256] NET05[257] 
+ NET05[258] NET05[259] NET05[260] NET05[261] NET05[262] NET05[263] NET05[264] 
+ NET05[265] NET05[266] NET05[267] NET05[268] NET05[269] NET05[270] NET05[271] 
+ NET05[272] NET05[273] NET05[274] NET05[275] NET05[276] NET05[277] NET05[278] 
+ NET05[279] NET05[280] NET05[281] NET05[282] NET05[283] NET05[284] NET05[285] 
+ NET05[286] NET05[287] NET05[288] NET05[289] NET05[290] NET05[291] NET05[292] 
+ NET05[293] NET05[294] NET05[295] NET05[296] NET05[297] NET05[298] NET05[299] 
+ NET05[300] NET05[301] NET05[302] NET05[303] NET05[304] NET05[305] NET05[306] 
+ NET05[307] NET05[308] NET05[309] NET05[310] NET05[311] NET05[312] NET05[313] 
+ NET05[314] NET05[315] NET05[316] NET05[317] NET05[318] NET05[319] NET05[320] 
+ NET05[321] NET05[322] NET05[323] NET05[324] NET05[325] NET05[326] NET05[327] 
+ NET05[328] NET05[329] NET05[330] NET05[331] NET05[332] NET05[333] NET05[334] 
+ NET05[335] NET05[336] NET05[337] NET05[338] NET05[339] NET05[340] NET05[341] 
+ NET05[342] NET05[343] NET05[344] NET05[345] NET05[346] NET05[347] NET05[348] 
+ NET05[349] NET05[350] NET05[351] NET05[352] NET05[353] NET05[354] NET05[355] 
+ NET05[356] NET05[357] NET05[358] NET05[359] NET05[360] NET05[361] NET05[362] 
+ NET05[363] NET05[364] NET05[365] NET05[366] NET05[367] NET05[368] NET05[369] 
+ NET05[370] NET05[371] NET05[372] NET05[373] NET05[374] NET05[375] NET05[376] 
+ NET05[377] NET05[378] NET05[379] NET05[380] NET05[381] NET05[382] NET05[383] 
+ NET05[384] NET05[385] NET05[386] NET05[387] NET05[388] NET05[389] NET05[390] 
+ NET05[391] NET05[392] NET05[393] NET05[394] NET05[395] NET05[396] NET05[397] 
+ NET05[398] NET05[399] NET05[400] NET05[401] NET05[402] NET05[403] NET05[404] 
+ NET05[405] NET05[406] NET05[407] NET05[408] NET05[409] NET05[410] NET05[411] 
+ NET05[412] NET05[413] NET05[414] NET05[415] NET05[416] NET05[417] NET05[418] 
+ NET05[419] NET05[420] NET05[421] NET05[422] NET05[423] NET05[424] NET05[425] 
+ NET05[426] NET05[427] NET05[428] NET05[429] NET05[430] NET05[431] NET05[432] 
+ NET05[433] NET05[434] NET05[435] NET05[436] NET05[437] NET05[438] NET05[439] 
+ NET05[440] NET05[441] NET05[442] NET05[443] NET05[444] NET05[445] NET05[446] 
+ NET05[447] NET05[448] NET05[449] NET05[450] NET05[451] NET05[452] NET05[453] 
+ NET05[454] NET05[455] NET05[456] NET05[457] NET05[458] NET05[459] NET05[460] 
+ NET05[461] NET05[462] NET05[463] NET05[464] NET05[465] NET05[466] NET05[467] 
+ NET05[468] NET05[469] NET05[470] NET05[471] NET05[472] NET05[473] NET05[474] 
+ NET05[475] NET05[476] NET05[477] NET05[478] NET05[479] NET05[480] NET05[481] 
+ NET05[482] NET05[483] NET05[484] NET05[485] NET05[486] NET05[487] NET05[488] 
+ NET05[489] NET05[490] NET05[491] NET05[492] NET05[493] NET05[494] NET05[495] 
+ NET05[496] NET05[497] NET05[498] NET05[499] NET05[500] NET05[501] NET05[502] 
+ NET05[503] NET05[504] NET05[505] NET05[506] NET05[507] NET05[508] NET05[509] 
+ NET05[510] NET05[511] NET07 NET011 S1AHSF400W40_TKBL_S384_CHAR
XI15 NET070 NET067 NET066 NET072[0] NET072[1] NET072[2] NET072[3] NET072[4] 
+ NET072[5] NET072[6] NET072[7] NET072[8] NET072[9] NET072[10] NET072[11] 
+ NET072[12] NET072[13] NET072[14] NET072[15] NET072[16] NET072[17] NET072[18] 
+ NET072[19] NET072[20] NET072[21] NET072[22] NET072[23] NET072[24] NET072[25] 
+ NET072[26] NET072[27] NET072[28] NET072[29] NET072[30] NET072[31] NET072[32] 
+ NET072[33] NET072[34] NET072[35] NET072[36] NET072[37] NET072[38] NET072[39] 
+ NET072[40] NET072[41] NET072[42] NET072[43] NET072[44] NET072[45] NET072[46] 
+ NET072[47] NET072[48] NET072[49] NET072[50] NET072[51] NET072[52] NET072[53] 
+ NET072[54] NET072[55] NET072[56] NET072[57] NET072[58] NET072[59] NET072[60] 
+ NET072[61] NET072[62] NET072[63] NET072[64] NET072[65] NET072[66] NET072[67] 
+ NET072[68] NET072[69] NET072[70] NET072[71] NET072[72] NET072[73] NET072[74] 
+ NET072[75] NET072[76] NET072[77] NET072[78] NET072[79] NET072[80] NET072[81] 
+ NET072[82] NET072[83] NET072[84] NET072[85] NET072[86] NET072[87] NET072[88] 
+ NET072[89] NET072[90] NET072[91] NET072[92] NET072[93] NET072[94] NET072[95] 
+ NET072[96] NET072[97] NET072[98] NET072[99] NET072[100] NET072[101] 
+ NET072[102] NET072[103] NET072[104] NET072[105] NET072[106] NET072[107] 
+ NET072[108] NET072[109] NET072[110] NET072[111] NET072[112] NET072[113] 
+ NET072[114] NET072[115] NET072[116] NET072[117] NET072[118] NET072[119] 
+ NET072[120] NET072[121] NET072[122] NET072[123] NET072[124] NET072[125] 
+ NET072[126] NET072[127] NET072[128] NET072[129] NET072[130] NET072[131] 
+ NET072[132] NET072[133] NET072[134] NET072[135] NET072[136] NET072[137] 
+ NET072[138] NET072[139] NET072[140] NET072[141] NET072[142] NET072[143] 
+ NET072[144] NET072[145] NET072[146] NET072[147] NET072[148] NET072[149] 
+ NET072[150] NET072[151] NET072[152] NET072[153] NET072[154] NET072[155] 
+ NET072[156] NET072[157] NET072[158] NET072[159] NET072[160] NET072[161] 
+ NET072[162] NET072[163] NET072[164] NET072[165] NET072[166] NET072[167] 
+ NET072[168] NET072[169] NET072[170] NET072[171] NET072[172] NET072[173] 
+ NET072[174] NET072[175] NET072[176] NET072[177] NET072[178] NET072[179] 
+ NET072[180] NET072[181] NET072[182] NET072[183] NET072[184] NET072[185] 
+ NET072[186] NET072[187] NET072[188] NET072[189] NET072[190] NET072[191] 
+ NET072[192] NET072[193] NET072[194] NET072[195] NET072[196] NET072[197] 
+ NET072[198] NET072[199] NET072[200] NET072[201] NET072[202] NET072[203] 
+ NET072[204] NET072[205] NET072[206] NET072[207] NET072[208] NET072[209] 
+ NET072[210] NET072[211] NET072[212] NET072[213] NET072[214] NET072[215] 
+ NET072[216] NET072[217] NET072[218] NET072[219] NET072[220] NET072[221] 
+ NET072[222] NET072[223] NET072[224] NET072[225] NET072[226] NET072[227] 
+ NET072[228] NET072[229] NET072[230] NET072[231] NET072[232] NET072[233] 
+ NET072[234] NET072[235] NET072[236] NET072[237] NET072[238] NET072[239] 
+ NET072[240] NET072[241] NET072[242] NET072[243] NET072[244] NET072[245] 
+ NET072[246] NET072[247] NET072[248] NET072[249] NET072[250] NET072[251] 
+ NET072[252] NET072[253] NET072[254] NET072[255] NET072[256] NET072[257] 
+ NET072[258] NET072[259] NET072[260] NET072[261] NET072[262] NET072[263] 
+ NET072[264] NET072[265] NET072[266] NET072[267] NET072[268] NET072[269] 
+ NET072[270] NET072[271] NET072[272] NET072[273] NET072[274] NET072[275] 
+ NET072[276] NET072[277] NET072[278] NET072[279] NET072[280] NET072[281] 
+ NET072[282] NET072[283] NET072[284] NET072[285] NET072[286] NET072[287] 
+ NET072[288] NET072[289] NET072[290] NET072[291] NET072[292] NET072[293] 
+ NET072[294] NET072[295] NET072[296] NET072[297] NET072[298] NET072[299] 
+ NET072[300] NET072[301] NET072[302] NET072[303] NET072[304] NET072[305] 
+ NET072[306] NET072[307] NET072[308] NET072[309] NET072[310] NET072[311] 
+ NET072[312] NET072[313] NET072[314] NET072[315] NET072[316] NET072[317] 
+ NET072[318] NET072[319] NET072[320] NET072[321] NET072[322] NET072[323] 
+ NET072[324] NET072[325] NET072[326] NET072[327] NET072[328] NET072[329] 
+ NET072[330] NET072[331] NET072[332] NET072[333] NET072[334] NET072[335] 
+ NET072[336] NET072[337] NET072[338] NET072[339] NET072[340] NET072[341] 
+ NET072[342] NET072[343] NET072[344] NET072[345] NET072[346] NET072[347] 
+ NET072[348] NET072[349] NET072[350] NET072[351] NET072[352] NET072[353] 
+ NET072[354] NET072[355] NET072[356] NET072[357] NET072[358] NET072[359] 
+ NET072[360] NET072[361] NET072[362] NET072[363] NET072[364] NET072[365] 
+ NET072[366] NET072[367] NET072[368] NET072[369] NET072[370] NET072[371] 
+ NET072[372] NET072[373] NET072[374] NET072[375] NET072[376] NET072[377] 
+ NET072[378] NET072[379] NET072[380] NET072[381] NET072[382] NET072[383] 
+ NET072[384] NET072[385] NET072[386] NET072[387] NET072[388] NET072[389] 
+ NET072[390] NET072[391] NET072[392] NET072[393] NET072[394] NET072[395] 
+ NET072[396] NET072[397] NET072[398] NET072[399] NET072[400] NET072[401] 
+ NET072[402] NET072[403] NET072[404] NET072[405] NET072[406] NET072[407] 
+ NET072[408] NET072[409] NET072[410] NET072[411] NET072[412] NET072[413] 
+ NET072[414] NET072[415] NET072[416] NET072[417] NET072[418] NET072[419] 
+ NET072[420] NET072[421] NET072[422] NET072[423] NET072[424] NET072[425] 
+ NET072[426] NET072[427] NET072[428] NET072[429] NET072[430] NET072[431] 
+ NET072[432] NET072[433] NET072[434] NET072[435] NET072[436] NET072[437] 
+ NET072[438] NET072[439] NET072[440] NET072[441] NET072[442] NET072[443] 
+ NET072[444] NET072[445] NET072[446] NET072[447] NET072[448] NET072[449] 
+ NET072[450] NET072[451] NET072[452] NET072[453] NET072[454] NET072[455] 
+ NET072[456] NET072[457] NET072[458] NET072[459] NET072[460] NET072[461] 
+ NET072[462] NET072[463] NET072[464] NET072[465] NET072[466] NET072[467] 
+ NET072[468] NET072[469] NET072[470] NET072[471] NET072[472] NET072[473] 
+ NET072[474] NET072[475] NET072[476] NET072[477] NET072[478] NET072[479] 
+ NET072[480] NET072[481] NET072[482] NET072[483] NET072[484] NET072[485] 
+ NET072[486] NET072[487] NET072[488] NET072[489] NET072[490] NET072[491] 
+ NET072[492] NET072[493] NET072[494] NET072[495] NET072[496] NET072[497] 
+ NET072[498] NET072[499] NET072[500] NET072[501] NET072[502] NET072[503] 
+ NET072[504] NET072[505] NET072[506] NET072[507] NET072[508] NET072[509] 
+ NET072[510] NET072[511] NET071[0] NET071[1] NET071[2] NET071[3] NET071[4] 
+ NET071[5] NET071[6] NET071[7] NET071[8] NET071[9] NET071[10] NET071[11] 
+ NET071[12] NET071[13] NET071[14] NET071[15] NET071[16] NET071[17] NET071[18] 
+ NET071[19] NET071[20] NET071[21] NET071[22] NET071[23] NET071[24] NET071[25] 
+ NET071[26] NET071[27] NET071[28] NET071[29] NET071[30] NET071[31] NET071[32] 
+ NET071[33] NET071[34] NET071[35] NET071[36] NET071[37] NET071[38] NET071[39] 
+ NET071[40] NET071[41] NET071[42] NET071[43] NET071[44] NET071[45] NET071[46] 
+ NET071[47] NET071[48] NET071[49] NET071[50] NET071[51] NET071[52] NET071[53] 
+ NET071[54] NET071[55] NET071[56] NET071[57] NET071[58] NET071[59] NET071[60] 
+ NET071[61] NET071[62] NET071[63] NET071[64] NET071[65] NET071[66] NET071[67] 
+ NET071[68] NET071[69] NET071[70] NET071[71] NET071[72] NET071[73] NET071[74] 
+ NET071[75] NET071[76] NET071[77] NET071[78] NET071[79] NET071[80] NET071[81] 
+ NET071[82] NET071[83] NET071[84] NET071[85] NET071[86] NET071[87] NET071[88] 
+ NET071[89] NET071[90] NET071[91] NET071[92] NET071[93] NET071[94] NET071[95] 
+ NET071[96] NET071[97] NET071[98] NET071[99] NET071[100] NET071[101] 
+ NET071[102] NET071[103] NET071[104] NET071[105] NET071[106] NET071[107] 
+ NET071[108] NET071[109] NET071[110] NET071[111] NET071[112] NET071[113] 
+ NET071[114] NET071[115] NET071[116] NET071[117] NET071[118] NET071[119] 
+ NET071[120] NET071[121] NET071[122] NET071[123] NET071[124] NET071[125] 
+ NET071[126] NET071[127] NET071[128] NET071[129] NET071[130] NET071[131] 
+ NET071[132] NET071[133] NET071[134] NET071[135] NET071[136] NET071[137] 
+ NET071[138] NET071[139] NET071[140] NET071[141] NET071[142] NET071[143] 
+ NET071[144] NET071[145] NET071[146] NET071[147] NET071[148] NET071[149] 
+ NET071[150] NET071[151] NET071[152] NET071[153] NET071[154] NET071[155] 
+ NET071[156] NET071[157] NET071[158] NET071[159] NET071[160] NET071[161] 
+ NET071[162] NET071[163] NET071[164] NET071[165] NET071[166] NET071[167] 
+ NET071[168] NET071[169] NET071[170] NET071[171] NET071[172] NET071[173] 
+ NET071[174] NET071[175] NET071[176] NET071[177] NET071[178] NET071[179] 
+ NET071[180] NET071[181] NET071[182] NET071[183] NET071[184] NET071[185] 
+ NET071[186] NET071[187] NET071[188] NET071[189] NET071[190] NET071[191] 
+ NET071[192] NET071[193] NET071[194] NET071[195] NET071[196] NET071[197] 
+ NET071[198] NET071[199] NET071[200] NET071[201] NET071[202] NET071[203] 
+ NET071[204] NET071[205] NET071[206] NET071[207] NET071[208] NET071[209] 
+ NET071[210] NET071[211] NET071[212] NET071[213] NET071[214] NET071[215] 
+ NET071[216] NET071[217] NET071[218] NET071[219] NET071[220] NET071[221] 
+ NET071[222] NET071[223] NET071[224] NET071[225] NET071[226] NET071[227] 
+ NET071[228] NET071[229] NET071[230] NET071[231] NET071[232] NET071[233] 
+ NET071[234] NET071[235] NET071[236] NET071[237] NET071[238] NET071[239] 
+ NET071[240] NET071[241] NET071[242] NET071[243] NET071[244] NET071[245] 
+ NET071[246] NET071[247] NET071[248] NET071[249] NET071[250] NET071[251] 
+ NET071[252] NET071[253] NET071[254] NET071[255] NET071[256] NET071[257] 
+ NET071[258] NET071[259] NET071[260] NET071[261] NET071[262] NET071[263] 
+ NET071[264] NET071[265] NET071[266] NET071[267] NET071[268] NET071[269] 
+ NET071[270] NET071[271] NET071[272] NET071[273] NET071[274] NET071[275] 
+ NET071[276] NET071[277] NET071[278] NET071[279] NET071[280] NET071[281] 
+ NET071[282] NET071[283] NET071[284] NET071[285] NET071[286] NET071[287] 
+ NET071[288] NET071[289] NET071[290] NET071[291] NET071[292] NET071[293] 
+ NET071[294] NET071[295] NET071[296] NET071[297] NET071[298] NET071[299] 
+ NET071[300] NET071[301] NET071[302] NET071[303] NET071[304] NET071[305] 
+ NET071[306] NET071[307] NET071[308] NET071[309] NET071[310] NET071[311] 
+ NET071[312] NET071[313] NET071[314] NET071[315] NET071[316] NET071[317] 
+ NET071[318] NET071[319] NET071[320] NET071[321] NET071[322] NET071[323] 
+ NET071[324] NET071[325] NET071[326] NET071[327] NET071[328] NET071[329] 
+ NET071[330] NET071[331] NET071[332] NET071[333] NET071[334] NET071[335] 
+ NET071[336] NET071[337] NET071[338] NET071[339] NET071[340] NET071[341] 
+ NET071[342] NET071[343] NET071[344] NET071[345] NET071[346] NET071[347] 
+ NET071[348] NET071[349] NET071[350] NET071[351] NET071[352] NET071[353] 
+ NET071[354] NET071[355] NET071[356] NET071[357] NET071[358] NET071[359] 
+ NET071[360] NET071[361] NET071[362] NET071[363] NET071[364] NET071[365] 
+ NET071[366] NET071[367] NET071[368] NET071[369] NET071[370] NET071[371] 
+ NET071[372] NET071[373] NET071[374] NET071[375] NET071[376] NET071[377] 
+ NET071[378] NET071[379] NET071[380] NET071[381] NET071[382] NET071[383] 
+ NET071[384] NET071[385] NET071[386] NET071[387] NET071[388] NET071[389] 
+ NET071[390] NET071[391] NET071[392] NET071[393] NET071[394] NET071[395] 
+ NET071[396] NET071[397] NET071[398] NET071[399] NET071[400] NET071[401] 
+ NET071[402] NET071[403] NET071[404] NET071[405] NET071[406] NET071[407] 
+ NET071[408] NET071[409] NET071[410] NET071[411] NET071[412] NET071[413] 
+ NET071[414] NET071[415] NET071[416] NET071[417] NET071[418] NET071[419] 
+ NET071[420] NET071[421] NET071[422] NET071[423] NET071[424] NET071[425] 
+ NET071[426] NET071[427] NET071[428] NET071[429] NET071[430] NET071[431] 
+ NET071[432] NET071[433] NET071[434] NET071[435] NET071[436] NET071[437] 
+ NET071[438] NET071[439] NET071[440] NET071[441] NET071[442] NET071[443] 
+ NET071[444] NET071[445] NET071[446] NET071[447] NET071[448] NET071[449] 
+ NET071[450] NET071[451] NET071[452] NET071[453] NET071[454] NET071[455] 
+ NET071[456] NET071[457] NET071[458] NET071[459] NET071[460] NET071[461] 
+ NET071[462] NET071[463] NET071[464] NET071[465] NET071[466] NET071[467] 
+ NET071[468] NET071[469] NET071[470] NET071[471] NET071[472] NET071[473] 
+ NET071[474] NET071[475] NET071[476] NET071[477] NET071[478] NET071[479] 
+ NET071[480] NET071[481] NET071[482] NET071[483] NET071[484] NET071[485] 
+ NET071[486] NET071[487] NET071[488] NET071[489] NET071[490] NET071[491] 
+ NET071[492] NET071[493] NET071[494] NET071[495] NET071[496] NET071[497] 
+ NET071[498] NET071[499] NET071[500] NET071[501] NET071[502] NET071[503] 
+ NET071[504] NET071[505] NET071[506] NET071[507] NET071[508] NET071[509] 
+ NET071[510] NET071[511] NET069 NET068 S1AHSF400W40_TKBL_S512_CHAR
XI11 NET026 NET023 NET022 NET013[0] NET013[1] NET013[2] NET013[3] NET013[4] 
+ NET013[5] NET013[6] NET013[7] NET013[8] NET013[9] NET013[10] NET013[11] 
+ NET013[12] NET013[13] NET013[14] NET013[15] NET013[16] NET013[17] NET013[18] 
+ NET013[19] NET013[20] NET013[21] NET013[22] NET013[23] NET013[24] NET013[25] 
+ NET013[26] NET013[27] NET013[28] NET013[29] NET013[30] NET013[31] NET013[32] 
+ NET013[33] NET013[34] NET013[35] NET013[36] NET013[37] NET013[38] NET013[39] 
+ NET013[40] NET013[41] NET013[42] NET013[43] NET013[44] NET013[45] NET013[46] 
+ NET013[47] NET013[48] NET013[49] NET013[50] NET013[51] NET013[52] NET013[53] 
+ NET013[54] NET013[55] NET013[56] NET013[57] NET013[58] NET013[59] NET013[60] 
+ NET013[61] NET013[62] NET013[63] NET010[0] NET010[1] NET010[2] NET010[3] 
+ NET010[4] NET010[5] NET010[6] NET010[7] NET010[8] NET010[9] NET010[10] 
+ NET010[11] NET010[12] NET010[13] NET010[14] NET010[15] NET010[16] NET010[17] 
+ NET010[18] NET010[19] NET010[20] NET010[21] NET010[22] NET010[23] NET010[24] 
+ NET010[25] NET010[26] NET010[27] NET010[28] NET010[29] NET010[30] NET010[31] 
+ NET010[32] NET010[33] NET010[34] NET010[35] NET010[36] NET010[37] NET010[38] 
+ NET010[39] NET010[40] NET010[41] NET010[42] NET010[43] NET010[44] NET010[45] 
+ NET010[46] NET010[47] NET010[48] NET010[49] NET010[50] NET010[51] NET010[52] 
+ NET010[53] NET010[54] NET010[55] NET010[56] NET010[57] NET010[58] NET010[59] 
+ NET010[60] NET010[61] NET010[62] NET010[63] NET025 NET024 S1AHSF400W40_TKBL_S64_CHAR
XTKBL_S256 NET20 NET18 NET017 NET21[0] NET21[1] NET21[2] NET21[3] NET21[4] 
+ NET21[5] NET21[6] NET21[7] NET21[8] NET21[9] NET21[10] NET21[11] NET21[12] 
+ NET21[13] NET21[14] NET21[15] NET21[16] NET21[17] NET21[18] NET21[19] 
+ NET21[20] NET21[21] NET21[22] NET21[23] NET21[24] NET21[25] NET21[26] 
+ NET21[27] NET21[28] NET21[29] NET21[30] NET21[31] NET21[32] NET21[33] 
+ NET21[34] NET21[35] NET21[36] NET21[37] NET21[38] NET21[39] NET21[40] 
+ NET21[41] NET21[42] NET21[43] NET21[44] NET21[45] NET21[46] NET21[47] 
+ NET21[48] NET21[49] NET21[50] NET21[51] NET21[52] NET21[53] NET21[54] 
+ NET21[55] NET21[56] NET21[57] NET21[58] NET21[59] NET21[60] NET21[61] 
+ NET21[62] NET21[63] NET21[64] NET21[65] NET21[66] NET21[67] NET21[68] 
+ NET21[69] NET21[70] NET21[71] NET21[72] NET21[73] NET21[74] NET21[75] 
+ NET21[76] NET21[77] NET21[78] NET21[79] NET21[80] NET21[81] NET21[82] 
+ NET21[83] NET21[84] NET21[85] NET21[86] NET21[87] NET21[88] NET21[89] 
+ NET21[90] NET21[91] NET21[92] NET21[93] NET21[94] NET21[95] NET21[96] 
+ NET21[97] NET21[98] NET21[99] NET21[100] NET21[101] NET21[102] NET21[103] 
+ NET21[104] NET21[105] NET21[106] NET21[107] NET21[108] NET21[109] NET21[110] 
+ NET21[111] NET21[112] NET21[113] NET21[114] NET21[115] NET21[116] NET21[117] 
+ NET21[118] NET21[119] NET21[120] NET21[121] NET21[122] NET21[123] NET21[124] 
+ NET21[125] NET21[126] NET21[127] NET21[128] NET21[129] NET21[130] NET21[131] 
+ NET21[132] NET21[133] NET21[134] NET21[135] NET21[136] NET21[137] NET21[138] 
+ NET21[139] NET21[140] NET21[141] NET21[142] NET21[143] NET21[144] NET21[145] 
+ NET21[146] NET21[147] NET21[148] NET21[149] NET21[150] NET21[151] NET21[152] 
+ NET21[153] NET21[154] NET21[155] NET21[156] NET21[157] NET21[158] NET21[159] 
+ NET21[160] NET21[161] NET21[162] NET21[163] NET21[164] NET21[165] NET21[166] 
+ NET21[167] NET21[168] NET21[169] NET21[170] NET21[171] NET21[172] NET21[173] 
+ NET21[174] NET21[175] NET21[176] NET21[177] NET21[178] NET21[179] NET21[180] 
+ NET21[181] NET21[182] NET21[183] NET21[184] NET21[185] NET21[186] NET21[187] 
+ NET21[188] NET21[189] NET21[190] NET21[191] NET21[192] NET21[193] NET21[194] 
+ NET21[195] NET21[196] NET21[197] NET21[198] NET21[199] NET21[200] NET21[201] 
+ NET21[202] NET21[203] NET21[204] NET21[205] NET21[206] NET21[207] NET21[208] 
+ NET21[209] NET21[210] NET21[211] NET21[212] NET21[213] NET21[214] NET21[215] 
+ NET21[216] NET21[217] NET21[218] NET21[219] NET21[220] NET21[221] NET21[222] 
+ NET21[223] NET21[224] NET21[225] NET21[226] NET21[227] NET21[228] NET21[229] 
+ NET21[230] NET21[231] NET21[232] NET21[233] NET21[234] NET21[235] NET21[236] 
+ NET21[237] NET21[238] NET21[239] NET21[240] NET21[241] NET21[242] NET21[243] 
+ NET21[244] NET21[245] NET21[246] NET21[247] NET21[248] NET21[249] NET21[250] 
+ NET21[251] NET21[252] NET21[253] NET21[254] NET21[255] NET15[0] NET15[1] 
+ NET15[2] NET15[3] NET15[4] NET15[5] NET15[6] NET15[7] NET15[8] NET15[9] 
+ NET15[10] NET15[11] NET15[12] NET15[13] NET15[14] NET15[15] NET15[16] 
+ NET15[17] NET15[18] NET15[19] NET15[20] NET15[21] NET15[22] NET15[23] 
+ NET15[24] NET15[25] NET15[26] NET15[27] NET15[28] NET15[29] NET15[30] 
+ NET15[31] NET15[32] NET15[33] NET15[34] NET15[35] NET15[36] NET15[37] 
+ NET15[38] NET15[39] NET15[40] NET15[41] NET15[42] NET15[43] NET15[44] 
+ NET15[45] NET15[46] NET15[47] NET15[48] NET15[49] NET15[50] NET15[51] 
+ NET15[52] NET15[53] NET15[54] NET15[55] NET15[56] NET15[57] NET15[58] 
+ NET15[59] NET15[60] NET15[61] NET15[62] NET15[63] NET15[64] NET15[65] 
+ NET15[66] NET15[67] NET15[68] NET15[69] NET15[70] NET15[71] NET15[72] 
+ NET15[73] NET15[74] NET15[75] NET15[76] NET15[77] NET15[78] NET15[79] 
+ NET15[80] NET15[81] NET15[82] NET15[83] NET15[84] NET15[85] NET15[86] 
+ NET15[87] NET15[88] NET15[89] NET15[90] NET15[91] NET15[92] NET15[93] 
+ NET15[94] NET15[95] NET15[96] NET15[97] NET15[98] NET15[99] NET15[100] 
+ NET15[101] NET15[102] NET15[103] NET15[104] NET15[105] NET15[106] NET15[107] 
+ NET15[108] NET15[109] NET15[110] NET15[111] NET15[112] NET15[113] NET15[114] 
+ NET15[115] NET15[116] NET15[117] NET15[118] NET15[119] NET15[120] NET15[121] 
+ NET15[122] NET15[123] NET15[124] NET15[125] NET15[126] NET15[127] NET15[128] 
+ NET15[129] NET15[130] NET15[131] NET15[132] NET15[133] NET15[134] NET15[135] 
+ NET15[136] NET15[137] NET15[138] NET15[139] NET15[140] NET15[141] NET15[142] 
+ NET15[143] NET15[144] NET15[145] NET15[146] NET15[147] NET15[148] NET15[149] 
+ NET15[150] NET15[151] NET15[152] NET15[153] NET15[154] NET15[155] NET15[156] 
+ NET15[157] NET15[158] NET15[159] NET15[160] NET15[161] NET15[162] NET15[163] 
+ NET15[164] NET15[165] NET15[166] NET15[167] NET15[168] NET15[169] NET15[170] 
+ NET15[171] NET15[172] NET15[173] NET15[174] NET15[175] NET15[176] NET15[177] 
+ NET15[178] NET15[179] NET15[180] NET15[181] NET15[182] NET15[183] NET15[184] 
+ NET15[185] NET15[186] NET15[187] NET15[188] NET15[189] NET15[190] NET15[191] 
+ NET15[192] NET15[193] NET15[194] NET15[195] NET15[196] NET15[197] NET15[198] 
+ NET15[199] NET15[200] NET15[201] NET15[202] NET15[203] NET15[204] NET15[205] 
+ NET15[206] NET15[207] NET15[208] NET15[209] NET15[210] NET15[211] NET15[212] 
+ NET15[213] NET15[214] NET15[215] NET15[216] NET15[217] NET15[218] NET15[219] 
+ NET15[220] NET15[221] NET15[222] NET15[223] NET15[224] NET15[225] NET15[226] 
+ NET15[227] NET15[228] NET15[229] NET15[230] NET15[231] NET15[232] NET15[233] 
+ NET15[234] NET15[235] NET15[236] NET15[237] NET15[238] NET15[239] NET15[240] 
+ NET15[241] NET15[242] NET15[243] NET15[244] NET15[245] NET15[246] NET15[247] 
+ NET15[248] NET15[249] NET15[250] NET15[251] NET15[252] NET15[253] NET15[254] 
+ NET15[255] NET19 NET16 S1AHSF400W40_TKBL_S256_CHAR
XI12 NET019 NET016 NET015 NET08[0] NET08[1] NET08[2] NET08[3] NET08[4] 
+ NET08[5] NET08[6] NET08[7] NET08[8] NET08[9] NET08[10] NET08[11] NET08[12] 
+ NET08[13] NET08[14] NET08[15] NET08[16] NET08[17] NET08[18] NET08[19] 
+ NET08[20] NET08[21] NET08[22] NET08[23] NET08[24] NET08[25] NET08[26] 
+ NET08[27] NET08[28] NET08[29] NET08[30] NET08[31] NET04[0] NET04[1] NET04[2] 
+ NET04[3] NET04[4] NET04[5] NET04[6] NET04[7] NET04[8] NET04[9] NET04[10] 
+ NET04[11] NET04[12] NET04[13] NET04[14] NET04[15] NET04[16] NET04[17] 
+ NET04[18] NET04[19] NET04[20] NET04[21] NET04[22] NET04[23] NET04[24] 
+ NET04[25] NET04[26] NET04[27] NET04[28] NET04[29] NET04[30] NET04[31] NET018 
+ NET01 S1AHSF400W40_TKBL_S32_CHAR
XI10 NET033 NET030 NET029 NET012[0] NET012[1] NET012[2] NET012[3] NET012[4] 
+ NET012[5] NET012[6] NET012[7] NET012[8] NET012[9] NET012[10] NET012[11] 
+ NET012[12] NET012[13] NET012[14] NET012[15] NET012[16] NET012[17] NET012[18] 
+ NET012[19] NET012[20] NET012[21] NET012[22] NET012[23] NET012[24] NET012[25] 
+ NET012[26] NET012[27] NET012[28] NET012[29] NET012[30] NET012[31] NET012[32] 
+ NET012[33] NET012[34] NET012[35] NET012[36] NET012[37] NET012[38] NET012[39] 
+ NET012[40] NET012[41] NET012[42] NET012[43] NET012[44] NET012[45] NET012[46] 
+ NET012[47] NET012[48] NET012[49] NET012[50] NET012[51] NET012[52] NET012[53] 
+ NET012[54] NET012[55] NET012[56] NET012[57] NET012[58] NET012[59] NET012[60] 
+ NET012[61] NET012[62] NET012[63] NET012[64] NET012[65] NET012[66] NET012[67] 
+ NET012[68] NET012[69] NET012[70] NET012[71] NET012[72] NET012[73] NET012[74] 
+ NET012[75] NET012[76] NET012[77] NET012[78] NET012[79] NET012[80] NET012[81] 
+ NET012[82] NET012[83] NET012[84] NET012[85] NET012[86] NET012[87] NET012[88] 
+ NET012[89] NET012[90] NET012[91] NET012[92] NET012[93] NET012[94] NET012[95] 
+ NET012[96] NET012[97] NET012[98] NET012[99] NET012[100] NET012[101] 
+ NET012[102] NET012[103] NET012[104] NET012[105] NET012[106] NET012[107] 
+ NET012[108] NET012[109] NET012[110] NET012[111] NET012[112] NET012[113] 
+ NET012[114] NET012[115] NET012[116] NET012[117] NET012[118] NET012[119] 
+ NET012[120] NET012[121] NET012[122] NET012[123] NET012[124] NET012[125] 
+ NET012[126] NET012[127] NET09[0] NET09[1] NET09[2] NET09[3] NET09[4] 
+ NET09[5] NET09[6] NET09[7] NET09[8] NET09[9] NET09[10] NET09[11] NET09[12] 
+ NET09[13] NET09[14] NET09[15] NET09[16] NET09[17] NET09[18] NET09[19] 
+ NET09[20] NET09[21] NET09[22] NET09[23] NET09[24] NET09[25] NET09[26] 
+ NET09[27] NET09[28] NET09[29] NET09[30] NET09[31] NET09[32] NET09[33] 
+ NET09[34] NET09[35] NET09[36] NET09[37] NET09[38] NET09[39] NET09[40] 
+ NET09[41] NET09[42] NET09[43] NET09[44] NET09[45] NET09[46] NET09[47] 
+ NET09[48] NET09[49] NET09[50] NET09[51] NET09[52] NET09[53] NET09[54] 
+ NET09[55] NET09[56] NET09[57] NET09[58] NET09[59] NET09[60] NET09[61] 
+ NET09[62] NET09[63] NET09[64] NET09[65] NET09[66] NET09[67] NET09[68] 
+ NET09[69] NET09[70] NET09[71] NET09[72] NET09[73] NET09[74] NET09[75] 
+ NET09[76] NET09[77] NET09[78] NET09[79] NET09[80] NET09[81] NET09[82] 
+ NET09[83] NET09[84] NET09[85] NET09[86] NET09[87] NET09[88] NET09[89] 
+ NET09[90] NET09[91] NET09[92] NET09[93] NET09[94] NET09[95] NET09[96] 
+ NET09[97] NET09[98] NET09[99] NET09[100] NET09[101] NET09[102] NET09[103] 
+ NET09[104] NET09[105] NET09[106] NET09[107] NET09[108] NET09[109] NET09[110] 
+ NET09[111] NET09[112] NET09[113] NET09[114] NET09[115] NET09[116] NET09[117] 
+ NET09[118] NET09[119] NET09[120] NET09[121] NET09[122] NET09[123] NET09[124] 
+ NET09[125] NET09[126] NET09[127] NET032 NET031 S1AHSF400W40_TKBL_S128_CHAR
XI14 NET035 NET020 NET014 NET049[0] NET049[1] NET049[2] NET049[3] NET049[4] 
+ NET049[5] NET049[6] NET049[7] NET049[8] NET049[9] NET049[10] NET049[11] 
+ NET049[12] NET049[13] NET049[14] NET049[15] NET048[0] NET048[1] NET048[2] 
+ NET048[3] NET048[4] NET048[5] NET048[6] NET048[7] NET048[8] NET048[9] 
+ NET048[10] NET048[11] NET048[12] NET048[13] NET048[14] NET048[15] NET036 
+ NET021 S1AHSF400W40_TKBL_S16_CHAR
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    TKBL_TRKPRE
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TKBL_TRKPRE PD TRKBL TRKWL VDDHD VDDI VSSI ZH ZL
*.PININFO PD:I TRKWL:I VDDHD:I ZH:O ZL:O TRKBL:B VDDI:B VSSI:B
MM0 ZH NET32 VDDI VDDI PCH L=60N W=6U M=1
MP0 TRKBL TRKWL VDDHD VDDI PCH L=60N W=3U M=1
MP1 NET28 NET28 VDDI VDDI PCH L=60N W=300N M=1
MP2 VDDI NET32 NET28 VDDI PCH L=60N W=300N M=1
MP3 NET14 NET17 VDDI VDDI PCH L=60N W=300N M=1
MN1 VSSI NET14 ZL VSSI NCH L=60N W=6U M=1
MM3 VSSI NET14 NET17 VSSI NCH L=60N W=300N M=1
MM2 NET17 NET17 VSSI VSSI NCH L=60N W=300N M=1
MM5 NET32 NET28 VSSI VSSI NCH L=60N W=300N M=1
MM1 TRKWL PD VSSI VSSI NCH L=60N W=300N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    TRKPRE_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TRKPRE_SIM PD TRKBL TRKWL VDDHD VDDI VSSI ZH ZL
*.PININFO PD:I TRKWL:I VDDHD:I ZH:O ZL:O TRKBL:B VDDI:B VSSI:B
XI1 NET23 TRKBL NET17 NET24 NET19 NET18 NET22 NET21 S1AHSF400W40_TKBL_TRKPRE
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    XDRV_STRAP_882_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_XDRV_STRAP_882_SB DEC_X2[0] DEC_X2_SHARE[0] VDDHD VDDI VSSI
*.PININFO DEC_X2[0]:B DEC_X2_SHARE[0]:B VDDHD:B VDDI:B VSSI:B
MM1 DEC_X2_SHARE[0] DEC_X2[0] VDDHD VDDI PCH L=60N W=4U M=2
MM10 DEC_X2_SHARE[0] DEC_X2[0] VSSI VSSI NCH L=60N W=4U M=2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    XDRV_LA512_882_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_XDRV_LA512_882_SB DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2_SHARE 
+ PD_BUF VDDHD VDDI VSSI WLOUT[0] WLOUT[1]
*.PININFO PD_BUF:I WLOUT[0]:O WLOUT[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B 
*.PININFO DEC_X0[3]:B DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B 
*.PININFO DEC_X1[0]:B DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B 
*.PININFO DEC_X1[5]:B DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B 
*.PININFO DEC_X2_SHARE:B VDDHD:B VDDI:B VSSI:B
MM0 VDDI DEC_X1[0] MWL0A VDDI PCH L=60N W=300N M=1
MM6 VDDI DEC_X1[0] MWL0 VDDI PCH L=60N W=300N M=1
MM3 VDDI DEC_X2[0] MWL0A VDDI PCH L=60N W=500N M=2
MM7 VDDI DEC_X0[0] MWL0 VDDI PCH L=60N W=300N M=1
MM1 WLOUT[1] MWL0A VDDHD VDDI PCH L=60N W=4U M=4
MP4 VDDHD PD_BUF VDDI VDDI PCH L=60N W=1U M=4
MM5 VDDI DEC_X0[1] MWL0A VDDI PCH L=60N W=300N M=1
MP19 VDDI DEC_X2[0] MWL0 VDDI PCH L=60N W=500N M=2
MM8 WLOUT[0] MWL0 VDDHD VDDI PCH L=60N W=4U M=4
MM2 WLOUT[1] MWL0A VSSI VSSI NCH L=60N W=4U M=2
MM11 SHARE DEC_X1[0] DEC_X2_SHARE VSSI NCH L=60N W=2U M=4
MN0 MWL0 DEC_X0[0] SHARE VSSI NCH L=60N W=4U M=1
MM9 WLOUT[0] MWL0 VSSI VSSI NCH L=60N W=4U M=2
MM4 MWL0A DEC_X0[1] SHARE VSSI NCH L=60N W=4U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_882_D
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_882_D DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2_SHARE 
+ PD_BUF VDDHD VDDI VSSI WL[0] WL[1]
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2_SHARE:B PD_BUF:B VDDHD:B 
*.PININFO VDDI:B VSSI:B WL[0]:B WL[1]:B
XSTRAP DEC_X2[0] DEC_X2_SHARE VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_882_SB
XWLDV DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI 
+ WL[0] WL[1] S1AHSF400W40_XDRV_LA512_882_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    XDRV_STRAP_884_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_XDRV_STRAP_884_SB DEC_X2[0] DEC_X2_SHARE[0] VDDHD VDDI VSSI
*.PININFO DEC_X2[0]:B DEC_X2_SHARE[0]:B VDDHD:B VDDI:B VSSI:B
MM1 DEC_X2_SHARE[0] DEC_X2[0] VDDHD VDDI PCH L=60N W=4U M=2
MM10 DEC_X2_SHARE[0] DEC_X2[0] VSSI VSSI NCH L=60N W=4U M=2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    XDRV_LA512_884_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_XDRV_LA512_884_SB DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WLOUT[0] WLOUT[1]
*.PININFO PD_BUF:I WLOUT[0]:O WLOUT[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B 
*.PININFO DEC_X0[3]:B DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B 
*.PININFO DEC_X1[0]:B DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B 
*.PININFO DEC_X1[5]:B DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B 
*.PININFO DEC_X2[2]:B DEC_X2[3]:B DEC_X2_SHARE:B VDDHD:B VDDI:B VSSI:B
MM9 WLOUT[0] MWL0 VSSI VSSI NCH L=60N W=4U M=2
MM11 SHARE DEC_X1[0] DEC_X2_SHARE VSSI NCH L=60N W=2U M=4
MM2 WLOUT[1] MWL0A VSSI VSSI NCH L=60N W=4U M=2
MM4 MWL0A DEC_X0[1] SHARE VSSI NCH L=60N W=4U M=1
MN0 MWL0 DEC_X0[0] SHARE VSSI NCH L=60N W=4U M=1
MM3 VDDI DEC_X2[0] MWL0A VDDI PCH L=60N W=500N M=2
MM1 WLOUT[1] MWL0A VDDHD VDDI PCH L=60N W=4U M=4
MM5 VDDI DEC_X0[1] MWL0A VDDI PCH L=60N W=300N M=1
MM6 VDDI DEC_X1[0] MWL0 VDDI PCH L=60N W=300N M=1
MM8 WLOUT[0] MWL0 VDDHD VDDI PCH L=60N W=4U M=4
MM0 VDDI DEC_X1[0] MWL0A VDDI PCH L=60N W=300N M=1
MM7 VDDI DEC_X0[0] MWL0 VDDI PCH L=60N W=300N M=1
MP4 VDDHD PD_BUF VDDI VDDI PCH L=60N W=1U M=4
MP19 VDDI DEC_X2[0] MWL0 VDDI PCH L=60N W=500N M=2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_884_D
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_884_D DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[0] WL[1]
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2_SHARE:B PD_BUF:B VDDHD:B VDDI:B VSSI:B WL[0]:B WL[1]:B
XSTRAP DEC_X2[0] DEC_X2_SHARE VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_884_SB
XWLDV DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2_SHARE 
+ PD_BUF VDDHD VDDI VSSI WL[0] WL[1] S1AHSF400W40_XDRV_LA512_884_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    XDRV_LA512_888_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_XDRV_LA512_888_SB DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_X2_SHARE PD_BUF VDDHD 
+ VDDI VSSI WLOUT[0] WLOUT[1]
*.PININFO PD_BUF:I WLOUT[0]:O WLOUT[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B 
*.PININFO DEC_X0[3]:B DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B 
*.PININFO DEC_X1[0]:B DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B 
*.PININFO DEC_X1[5]:B DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B 
*.PININFO DEC_X2[2]:B DEC_X2[3]:B DEC_X2[4]:B DEC_X2[5]:B DEC_X2[6]:B 
*.PININFO DEC_X2[7]:B DEC_X2_SHARE:B VDDHD:B VDDI:B VSSI:B
MM3 VDDI DEC_X2[0] MWL0A VDDI PCH L=60N W=500N M=2
MM0 VDDI DEC_X1[0] MWL0A VDDI PCH L=60N W=300N M=1
MM5 VDDI DEC_X0[1] MWL0A VDDI PCH L=60N W=300N M=1
MM6 VDDI DEC_X1[0] MWL0 VDDI PCH L=60N W=300N M=1
MP19 VDDI DEC_X2[0] MWL0 VDDI PCH L=60N W=500N M=2
MM1 WLOUT[1] MWL0A VDDHD VDDI PCH L=60N W=4U M=4
MP4 VDDHD PD_BUF VDDI VDDI PCH L=60N W=1U M=4
MM7 VDDI DEC_X0[0] MWL0 VDDI PCH L=60N W=300N M=1
MM8 WLOUT[0] MWL0 VDDHD VDDI PCH L=60N W=4U M=4
MM4 MWL0A DEC_X0[1] SHARE VSSI NCH L=60N W=4U M=1
MM2 WLOUT[1] MWL0A VSSI VSSI NCH L=60N W=4U M=2
MM11 SHARE DEC_X1[0] DEC_X2_SHARE VSSI NCH L=60N W=4U M=2
MM9 WLOUT[0] MWL0 VSSI VSSI NCH L=60N W=4U M=2
MN0 MWL0 DEC_X0[0] SHARE VSSI NCH L=60N W=4U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    XDRV_STRAP_888_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_XDRV_STRAP_888_SB DEC_X2[0] DEC_X2_SHARE[0] VDDHD VDDI VSSI
*.PININFO DEC_X2[0]:B DEC_X2_SHARE[0]:B VDDHD:B VDDI:B VSSI:B
MM1 DEC_X2_SHARE[0] DEC_X2[0] VDDHD VDDI PCH L=60N W=4U M=2
MM3 DEC_X2_SHARE[0] DEC_X2[0] VSSI VSSI NCH L=60N W=1U M=2
MM10 DEC_X2_SHARE[0] DEC_X2[0] VSSI VSSI NCH L=60N W=4U M=2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_888_D
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_888_D DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_X2_SHARE PD_BUF VDDHD 
+ VDDI VSSI WL[0] WL[1]
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2[4]:B DEC_X2[5]:B DEC_X2[6]:B DEC_X2[7]:B DEC_X2_SHARE:B 
*.PININFO PD_BUF:B VDDHD:B VDDI:B VSSI:B WL[0]:B WL[1]:B
XWLDV DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] 
+ DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[0] 
+ WL[1] S1AHSF400W40_XDRV_LA512_888_SB
XSTRAP DEC_X2[0] DEC_X2_SHARE VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_888_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_D_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_D_SIM DEC_X0_BT[0] DEC_X0_BT[1] DEC_X0_BT[2] DEC_X0_BT[3] 
+ DEC_X0_BT[4] DEC_X0_BT[5] DEC_X0_BT[6] DEC_X0_BT[7] DEC_X0_TP[0] 
+ DEC_X0_TP[1] DEC_X0_TP[2] DEC_X0_TP[3] DEC_X0_TP[4] DEC_X0_TP[5] 
+ DEC_X0_TP[6] DEC_X0_TP[7] DEC_X1_BT[0] DEC_X1_BT[1] DEC_X1_BT[2] 
+ DEC_X1_BT[3] DEC_X1_BT[4] DEC_X1_BT[5] DEC_X1_BT[6] DEC_X1_BT[7] 
+ DEC_X1_TP[0] DEC_X1_TP[1] DEC_X1_TP[2] DEC_X1_TP[3] DEC_X1_TP[4] 
+ DEC_X1_TP[5] DEC_X1_TP[6] DEC_X1_TP[7] DEC_X2_BT[0] DEC_X2_BT[1] 
+ DEC_X2_BT[2] DEC_X2_BT[3] DEC_X2_BT[4] DEC_X2_BT[5] DEC_X2_BT[6] 
+ DEC_X2_BT[7] DEC_X2_SHARE_TP DEC_X2_TP[0] DEC_X2_TP[1] DEC_X2_TP[2] 
+ DEC_X2_TP[3] DEC_X2_TP[4] DEC_X2_TP[5] DEC_X2_TP[6] DEC_X2_TP[7] PD_BUF_BT 
+ PD_BUF_TP VDDHD VDDI VSSI WL_LT[0] WL_LT[1] WL_RT[0] WL_RT[1]
*.PININFO DEC_X0_BT[0]:I DEC_X0_BT[1]:I DEC_X0_BT[2]:I DEC_X0_BT[3]:I 
*.PININFO DEC_X0_BT[4]:I DEC_X0_BT[5]:I DEC_X0_BT[6]:I DEC_X0_BT[7]:I 
*.PININFO DEC_X1_BT[0]:I DEC_X1_BT[1]:I DEC_X1_BT[2]:I DEC_X1_BT[3]:I 
*.PININFO DEC_X1_BT[4]:I DEC_X1_BT[5]:I DEC_X1_BT[6]:I DEC_X1_BT[7]:I 
*.PININFO PD_BUF_BT:I DEC_X0_TP[0]:O DEC_X0_TP[1]:O DEC_X0_TP[2]:O 
*.PININFO DEC_X0_TP[3]:O DEC_X0_TP[4]:O DEC_X0_TP[5]:O DEC_X0_TP[6]:O 
*.PININFO DEC_X0_TP[7]:O DEC_X1_TP[0]:O DEC_X1_TP[1]:O DEC_X1_TP[2]:O 
*.PININFO DEC_X1_TP[3]:O DEC_X1_TP[4]:O DEC_X1_TP[5]:O DEC_X1_TP[6]:O 
*.PININFO DEC_X1_TP[7]:O PD_BUF_TP:O DEC_X2_BT[0]:B DEC_X2_BT[1]:B 
*.PININFO DEC_X2_BT[2]:B DEC_X2_BT[3]:B DEC_X2_BT[4]:B DEC_X2_BT[5]:B 
*.PININFO DEC_X2_BT[6]:B DEC_X2_BT[7]:B DEC_X2_SHARE_TP:B DEC_X2_TP[0]:B 
*.PININFO DEC_X2_TP[1]:B DEC_X2_TP[2]:B DEC_X2_TP[3]:B DEC_X2_TP[4]:B 
*.PININFO DEC_X2_TP[5]:B DEC_X2_TP[6]:B DEC_X2_TP[7]:B VDDHD:B VDDI:B VSSI:B 
*.PININFO WL_LT[0]:B WL_LT[1]:B WL_RT[0]:B WL_RT[1]:B
XI26 NET025[0] NET025[1] NET025[2] NET025[3] NET025[4] NET025[5] NET025[6] 
+ NET025[7] NET030[0] NET030[1] NET030[2] NET030[3] NET030[4] NET030[5] 
+ NET030[6] NET030[7] NET027[0] NET027[1] NET026 NET01 NET08 NET02 NET06 
+ NET07[0] NET07[1] S1AHSF400W40_SB_WLDV_882_D
XI25 NET04[0] NET04[1] NET04[2] NET04[3] NET04[4] NET04[5] NET04[6] NET04[7] 
+ NET05[0] NET05[1] NET05[2] NET05[3] NET05[4] NET05[5] NET05[6] NET05[7] 
+ NET010[0] NET010[1] NET010[2] NET010[3] NET03 NET018 NET023 NET022 NET021 
+ NET019[0] NET019[1] S1AHSF400W40_SB_WLDV_884_D
XI27 NET045[0] NET045[1] NET045[2] NET045[3] NET045[4] NET045[5] NET045[6] 
+ NET045[7] NET043[0] NET043[1] NET043[2] NET043[3] NET043[4] NET043[5] 
+ NET043[6] NET043[7] NET044[0] NET044[1] NET044[2] NET044[3] NET044[4] 
+ NET044[5] NET044[6] NET044[7] NET046 NET038 NET042 NET041 NET040 NET039[0] 
+ NET039[1] S1AHSF400W40_SB_WLDV_888_D
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_882_U_64
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_882_U_64 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2_SHARE 
+ PD_BUF VDDHD VDDI VSSI WL[0] WL[1]
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2_SHARE:B PD_BUF:B VDDHD:B 
*.PININFO VDDI:B VSSI:B WL[0]:B WL[1]:B
XWLDV DEC_X0[6] DEC_X0[7] NET15[0] NET15[1] NET15[2] NET15[3] NET15[4] 
+ NET15[5] DEC_X1[7] NET12[0] NET12[1] NET12[2] NET12[3] NET12[4] NET12[5] 
+ NET12[6] DEC_X2[0] NET10 DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[0] WL[1] 
+ S1AHSF400W40_XDRV_LA512_882_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_882_U_66
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_882_U_66 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2_SHARE 
+ PD_BUF VDDHD VDDI VSSI WL[0] WL[1]
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2_SHARE:B PD_BUF:B VDDHD:B 
*.PININFO VDDI:B VSSI:B WL[0]:B WL[1]:B
XWLDV DEC_X0[0] DEC_X0[1] NET15[0] NET15[1] NET15[2] NET15[3] NET15[4] 
+ NET15[5] DEC_X1[0] NET12[0] NET12[1] NET12[2] NET12[3] NET12[4] NET12[5] 
+ NET12[6] DEC_X2[1] NET10 DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[0] WL[1] 
+ S1AHSF400W40_XDRV_LA512_882_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_888_U_384
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_888_U_384 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_X2_SHARE PD_BUF VDDHD 
+ VDDI VSSI WL[0] WL[1]
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2[4]:B DEC_X2[5]:B DEC_X2[6]:B DEC_X2[7]:B DEC_X2_SHARE:B 
*.PININFO PD_BUF:B VDDHD:B VDDI:B VSSI:B WL[0]:B WL[1]:B
XWLDV DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X2[5] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ DEC_X2[4] DEC_X2[6] DEC_X2[7] DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[0] 
+ WL[1] S1AHSF400W40_XDRV_LA512_888_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_888_U_386
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_888_U_386 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_X2_SHARE PD_BUF VDDHD 
+ VDDI VSSI WL[0] WL[1]
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2[4]:B DEC_X2[5]:B DEC_X2[6]:B DEC_X2[7]:B DEC_X2_SHARE:B 
*.PININFO PD_BUF:B VDDHD:B VDDI:B VSSI:B WL[0]:B WL[1]:B
XWLDV DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ DEC_X2[4] DEC_X2[5] DEC_X2[7] DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[0] 
+ WL[1] S1AHSF400W40_XDRV_LA512_888_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_882_U_128
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_882_U_128 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2_SHARE 
+ PD_BUF VDDHD VDDI VSSI WL[0] WL[1]
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2_SHARE:B PD_BUF:B VDDHD:B 
*.PININFO VDDI:B VSSI:B WL[0]:B WL[1]:B
XWLDV DEC_X0[6] DEC_X0[7] NET15[0] NET15[1] NET15[2] NET15[3] NET15[4] 
+ NET15[5] DEC_X1[7] NET12[0] NET12[1] NET12[2] NET12[3] NET12[4] NET12[5] 
+ NET12[6] DEC_X2[1] NET10 DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[0] WL[1] 
+ S1AHSF400W40_XDRV_LA512_882_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_882_U_16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_882_U_16 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2_SHARE 
+ PD_BUF VDDHD VDDI VSSI WL[0] WL[1]
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2_SHARE:B PD_BUF:B VDDHD:B 
*.PININFO VDDI:B VSSI:B WL[0]:B WL[1]:B
XWLDV DEC_X0[6] DEC_X0[7] NET15[0] NET15[1] NET15[2] NET15[3] NET15[4] 
+ NET15[5] DEC_X1[1] NET12[0] NET12[1] NET12[2] NET12[3] NET12[4] NET12[5] 
+ NET12[6] DEC_X2[0] NET10 DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[0] WL[1] 
+ S1AHSF400W40_XDRV_LA512_882_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_884_U_130
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_884_U_130 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[0] WL[1]
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2_SHARE:B PD_BUF:B VDDHD:B VDDI:B VSSI:B WL[0]:B WL[1]:B
XWLDV DEC_X0[0] DEC_X0[1] NET11[0] NET11[1] NET11[2] NET11[3] NET11[4] 
+ NET11[5] DEC_X1[0] NET13[0] NET13[1] NET13[2] NET13[3] NET13[4] NET13[5] 
+ NET13[6] DEC_X2[2] NET12[0] NET12[1] NET12[2] DEC_X2_SHARE PD_BUF VDDHD VDDI 
+ VSSI WL[0] WL[1] S1AHSF400W40_XDRV_LA512_884_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_884_U_256
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_884_U_256 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[0] WL[1]
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2_SHARE:B PD_BUF:B VDDHD:B VDDI:B VSSI:B WL[0]:B WL[1]:B
XWLDV DEC_X0[6] DEC_X0[7] NET11[0] NET11[1] NET11[2] NET11[3] NET11[4] 
+ NET11[5] DEC_X1[7] NET13[0] NET13[1] NET13[2] NET13[3] NET13[4] NET13[5] 
+ NET13[6] DEC_X2[3] NET12[0] NET12[1] NET12[2] DEC_X2_SHARE PD_BUF VDDHD VDDI 
+ VSSI WL[0] WL[1] S1AHSF400W40_XDRV_LA512_884_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_888_U_258
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_888_U_258 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_X2_SHARE PD_BUF VDDHD 
+ VDDI VSSI WL[0] WL[1]
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2[4]:B DEC_X2[5]:B DEC_X2[6]:B DEC_X2[7]:B DEC_X2_SHARE:B 
*.PININFO PD_BUF:B VDDHD:B VDDI:B VSSI:B WL[0]:B WL[1]:B
XWLDV DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[4] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[0] 
+ WL[1] S1AHSF400W40_XDRV_LA512_888_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_888_U_512
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_888_U_512 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_X2_SHARE PD_BUF VDDHD 
+ VDDI VSSI WL[0] WL[1]
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2[4]:B DEC_X2[5]:B DEC_X2[6]:B DEC_X2[7]:B DEC_X2_SHARE:B 
*.PININFO PD_BUF:B VDDHD:B VDDI:B VSSI:B WL[0]:B WL[1]:B
XWLDV DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X2[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[0] 
+ WL[1] S1AHSF400W40_XDRV_LA512_888_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_U_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_U_SIM DEC_X0_BT[0] DEC_X0_BT[1] DEC_X0_BT[2] DEC_X0_BT[3] 
+ DEC_X0_BT[4] DEC_X0_BT[5] DEC_X0_BT[6] DEC_X0_BT[7] DEC_X0_TP[0] 
+ DEC_X0_TP[1] DEC_X0_TP[2] DEC_X0_TP[3] DEC_X0_TP[4] DEC_X0_TP[5] 
+ DEC_X0_TP[6] DEC_X0_TP[7] DEC_X1_BT[0] DEC_X1_BT[1] DEC_X1_BT[2] 
+ DEC_X1_BT[3] DEC_X1_BT[4] DEC_X1_BT[5] DEC_X1_BT[6] DEC_X1_BT[7] 
+ DEC_X1_TP[0] DEC_X1_TP[1] DEC_X1_TP[2] DEC_X1_TP[3] DEC_X1_TP[4] 
+ DEC_X1_TP[5] DEC_X1_TP[6] DEC_X1_TP[7] DEC_X2_BT[0] DEC_X2_BT[1] 
+ DEC_X2_BT[2] DEC_X2_BT[3] DEC_X2_BT[4] DEC_X2_BT[5] DEC_X2_BT[6] 
+ DEC_X2_BT[7] DEC_X2_SHARE_BT DEC_X2_SHARE_TP DEC_X2_TP[0] DEC_X2_TP[1] 
+ DEC_X2_TP[2] DEC_X2_TP[3] DEC_X2_TP[4] DEC_X2_TP[5] DEC_X2_TP[6] 
+ DEC_X2_TP[7] PD_BUF_BT PD_BUF_TP VDDHD VDDI VSSI WL_LT[0] WL_LT[1] WL_RT[0] 
+ WL_RT[1]
*.PININFO DEC_X0_BT[0]:I DEC_X0_BT[1]:I DEC_X0_BT[2]:I DEC_X0_BT[3]:I 
*.PININFO DEC_X0_BT[4]:I DEC_X0_BT[5]:I DEC_X0_BT[6]:I DEC_X0_BT[7]:I 
*.PININFO DEC_X1_BT[0]:I DEC_X1_BT[1]:I DEC_X1_BT[2]:I DEC_X1_BT[3]:I 
*.PININFO DEC_X1_BT[4]:I DEC_X1_BT[5]:I DEC_X1_BT[6]:I DEC_X1_BT[7]:I 
*.PININFO PD_BUF_BT:I DEC_X0_TP[0]:O DEC_X0_TP[1]:O DEC_X0_TP[2]:O 
*.PININFO DEC_X0_TP[3]:O DEC_X0_TP[4]:O DEC_X0_TP[5]:O DEC_X0_TP[6]:O 
*.PININFO DEC_X0_TP[7]:O DEC_X1_TP[0]:O DEC_X1_TP[1]:O DEC_X1_TP[2]:O 
*.PININFO DEC_X1_TP[3]:O DEC_X1_TP[4]:O DEC_X1_TP[5]:O DEC_X1_TP[6]:O 
*.PININFO DEC_X1_TP[7]:O PD_BUF_TP:O DEC_X2_BT[0]:B DEC_X2_BT[1]:B 
*.PININFO DEC_X2_BT[2]:B DEC_X2_BT[3]:B DEC_X2_BT[4]:B DEC_X2_BT[5]:B 
*.PININFO DEC_X2_BT[6]:B DEC_X2_BT[7]:B DEC_X2_SHARE_BT:B DEC_X2_SHARE_TP:B 
*.PININFO DEC_X2_TP[0]:B DEC_X2_TP[1]:B DEC_X2_TP[2]:B DEC_X2_TP[3]:B 
*.PININFO DEC_X2_TP[4]:B DEC_X2_TP[5]:B DEC_X2_TP[6]:B DEC_X2_TP[7]:B VDDHD:B 
*.PININFO VDDI:B VSSI:B WL_LT[0]:B WL_LT[1]:B WL_RT[0]:B WL_RT[1]:B
XI36 NET011[0] NET011[1] NET011[2] NET011[3] NET011[4] NET011[5] NET011[6] 
+ NET011[7] NET055[0] NET055[1] NET055[2] NET055[3] NET055[4] NET055[5] 
+ NET055[6] NET055[7] NET08[0] NET08[1] NET051 NET013 NET010 NET025 NET05 
+ NET02[0] NET02[1] S1AHSF400W40_SB_WLDV_882_U_64
XI38 NET093[0] NET093[1] NET093[2] NET093[3] NET093[4] NET093[5] NET093[6] 
+ NET093[7] NET094[0] NET094[1] NET094[2] NET094[3] NET094[4] NET094[5] 
+ NET094[6] NET094[7] NET092[0] NET092[1] NET095 NET087 NET091 NET090 NET03 
+ NET06[0] NET06[1] S1AHSF400W40_SB_WLDV_882_U_66
XI40 NET0103[0] NET0103[1] NET0103[2] NET0103[3] NET0103[4] NET0103[5] 
+ NET0103[6] NET0103[7] NET0101[0] NET0101[1] NET0101[2] NET0101[3] NET0101[4] 
+ NET0101[5] NET0101[6] NET0101[7] NET0102[0] NET0102[1] NET0102[2] NET0102[3] 
+ NET0102[4] NET0102[5] NET0102[6] NET0102[7] NET0104 NET096 NET0100 NET099 
+ NET098 NET097[0] NET097[1] S1AHSF400W40_SB_WLDV_888_U_384
XI41 NET0112[0] NET0112[1] NET0112[2] NET0112[3] NET0112[4] NET0112[5] 
+ NET0112[6] NET0112[7] NET0110[0] NET0110[1] NET0110[2] NET0110[3] NET0110[4] 
+ NET0110[5] NET0110[6] NET0110[7] NET0111[0] NET0111[1] NET0111[2] NET0111[3] 
+ NET0111[4] NET0111[5] NET0111[6] NET0111[7] NET0113 NET0105 NET0109 NET0108 
+ NET0107 NET0106[0] NET0106[1] S1AHSF400W40_SB_WLDV_888_U_386
XI39 NET0120[0] NET0120[1] NET0120[2] NET0120[3] NET0120[4] NET0120[5] 
+ NET0120[6] NET0120[7] NET0121[0] NET0121[1] NET0121[2] NET0121[3] NET0121[4] 
+ NET0121[5] NET0121[6] NET0121[7] NET0119[0] NET0119[1] NET0122 NET0114 
+ NET0118 NET0117 NET0116 NET0115[0] NET0115[1] S1AHSF400W40_SB_WLDV_882_U_128
XI35 NET052[0] NET052[1] NET052[2] NET052[3] NET052[4] NET052[5] NET052[6] 
+ NET052[7] NET089[0] NET089[1] NET089[2] NET089[3] NET089[4] NET089[5] 
+ NET089[6] NET089[7] NET088[0] NET088[1] NET04 NET028 NET032 NET031 NET030 
+ NET029[0] NET029[1] S1AHSF400W40_SB_WLDV_882_U_16
XI32 NET022[0] NET022[1] NET022[2] NET022[3] NET022[4] NET022[5] NET022[6] 
+ NET022[7] NET021[0] NET021[1] NET021[2] NET021[3] NET021[4] NET021[5] 
+ NET021[6] NET021[7] NET01[0] NET01[1] NET01[2] NET01[3] NET023 NET016 NET020 
+ NET019 NET018 NET017[0] NET017[1] S1AHSF400W40_SB_WLDV_884_U_130
XI29 NET29[0] NET29[1] NET29[2] NET29[3] NET29[4] NET29[5] NET29[6] NET29[7] 
+ NET28[0] NET28[1] NET28[2] NET28[3] NET28[4] NET28[5] NET28[6] NET28[7] 
+ NET024[0] NET024[1] NET024[2] NET024[3] NET015 NET22 NET26 NET25 NET24 
+ NET014[0] NET014[1] S1AHSF400W40_SB_WLDV_884_U_256
XI33 NET040[0] NET040[1] NET040[2] NET040[3] NET040[4] NET040[5] NET040[6] 
+ NET040[7] NET038[0] NET038[1] NET038[2] NET038[3] NET038[4] NET038[5] 
+ NET038[6] NET038[7] NET039[0] NET039[1] NET039[2] NET039[3] NET039[4] 
+ NET039[5] NET039[6] NET039[7] NET041 NET033 NET037 NET036 NET035 NET034[0] 
+ NET034[1] S1AHSF400W40_SB_WLDV_888_U_258
XI34 NET049[0] NET049[1] NET049[2] NET049[3] NET049[4] NET049[5] NET049[6] 
+ NET049[7] NET047[0] NET047[1] NET047[2] NET047[3] NET047[4] NET047[5] 
+ NET047[6] NET047[7] NET048[0] NET048[1] NET048[2] NET048[3] NET048[4] 
+ NET048[5] NET048[6] NET048[7] NET050 NET042 NET046 NET045 NET044 NET043[0] 
+ NET043[1] S1AHSF400W40_SB_WLDV_888_U_512
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    XDRV_882_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_XDRV_882_SB DEC_X0[0] DEC_X0[1] DEC_X1 DEC_X2 DEC_X2_SHARE PD_BUF 
+ VDDHD VDDI VSSI WLOUT[0] WLOUT[1]
*.PININFO DEC_X0[0]:I DEC_X0[1]:I DEC_X1:I DEC_X2:I DEC_X2_SHARE:I PD_BUF:I 
*.PININFO WLOUT[0]:O WLOUT[1]:O VDDHD:B VDDI:B VSSI:B
XWLDV DEC_X0[0] DEC_X0[1] NET22[0] NET22[1] NET22[2] NET22[3] NET22[4] 
+ NET22[5] DEC_X1 NET18[0] NET18[1] NET18[2] NET18[3] NET18[4] NET18[5] 
+ NET18[6] DEC_X2 NET018 DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WLOUT[0] WLOUT[1] 
+ S1AHSF400W40_XDRV_LA512_882_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    WLDV_2X1_882_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_WLDV_2X1_882_SB DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1 DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[0] WL[1] WL[2] WL[3]
*.PININFO DEC_X0[0]:I DEC_X0[1]:I DEC_X0[2]:I DEC_X0[3]:I DEC_X1:I DEC_X2:I 
*.PININFO DEC_X2_SHARE:I PD_BUF:I WL[0]:O WL[1]:O WL[2]:O WL[3]:O VDDHD:B 
*.PININFO VDDI:B VSSI:B
XWLDV_0 DEC_X0[0] DEC_X0[1] DEC_X1 DEC_X2 DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI 
+ WL[0] WL[1] S1AHSF400W40_XDRV_882_SB
XWLDV_1 DEC_X0[2] DEC_X0[3] DEC_X1 DEC_X2 DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI 
+ WL[2] WL[3] S1AHSF400W40_XDRV_882_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    WLDV_64X1_882_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_WLDV_64X1_882_SB DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2 DEC_X2_SHARE PD_BUF VDDHD 
+ VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] 
+ WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] 
+ WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] 
+ WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] 
+ WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] 
+ WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63]
*.PININFO DEC_X0[0]:I DEC_X0[1]:I DEC_X0[2]:I DEC_X0[3]:I DEC_X0[4]:I 
*.PININFO DEC_X0[5]:I DEC_X0[6]:I DEC_X0[7]:I DEC_X1[0]:I DEC_X1[1]:I 
*.PININFO DEC_X1[2]:I DEC_X1[3]:I DEC_X1[4]:I DEC_X1[5]:I DEC_X1[6]:I 
*.PININFO DEC_X1[7]:I DEC_X2:I DEC_X2_SHARE:I PD_BUF:I WL[0]:O WL[1]:O WL[2]:O 
*.PININFO WL[3]:O WL[4]:O WL[5]:O WL[6]:O WL[7]:O WL[8]:O WL[9]:O WL[10]:O 
*.PININFO WL[11]:O WL[12]:O WL[13]:O WL[14]:O WL[15]:O WL[16]:O WL[17]:O 
*.PININFO WL[18]:O WL[19]:O WL[20]:O WL[21]:O WL[22]:O WL[23]:O WL[24]:O 
*.PININFO WL[25]:O WL[26]:O WL[27]:O WL[28]:O WL[29]:O WL[30]:O WL[31]:O 
*.PININFO WL[32]:O WL[33]:O WL[34]:O WL[35]:O WL[36]:O WL[37]:O WL[38]:O 
*.PININFO WL[39]:O WL[40]:O WL[41]:O WL[42]:O WL[43]:O WL[44]:O WL[45]:O 
*.PININFO WL[46]:O WL[47]:O WL[48]:O WL[49]:O WL[50]:O WL[51]:O WL[52]:O 
*.PININFO WL[53]:O WL[54]:O WL[55]:O WL[56]:O WL[57]:O WL[58]:O WL[59]:O 
*.PININFO WL[60]:O WL[61]:O WL[62]:O WL[63]:O VDDHD:B VDDI:B VSSI:B
XWLDV_2X1<0> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[0] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[0] WL[1] WL[2] WL[3] S1AHSF400W40_WLDV_2X1_882_SB
XWLDV_2X1<1> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[4] WL[5] WL[6] WL[7] S1AHSF400W40_WLDV_2X1_882_SB
XWLDV_2X1<2> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[1] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[8] WL[9] WL[10] WL[11] 
+ S1AHSF400W40_WLDV_2X1_882_SB
XWLDV_2X1<3> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[12] WL[13] WL[14] WL[15] 
+ S1AHSF400W40_WLDV_2X1_882_SB
XWLDV_2X1<4> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[2] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[16] WL[17] WL[18] WL[19] 
+ S1AHSF400W40_WLDV_2X1_882_SB
XWLDV_2X1<5> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[20] WL[21] WL[22] WL[23] 
+ S1AHSF400W40_WLDV_2X1_882_SB
XWLDV_2X1<6> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[3] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[24] WL[25] WL[26] WL[27] 
+ S1AHSF400W40_WLDV_2X1_882_SB
XWLDV_2X1<7> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[28] WL[29] WL[30] WL[31] 
+ S1AHSF400W40_WLDV_2X1_882_SB
XWLDV_2X1<8> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[4] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[32] WL[33] WL[34] WL[35] 
+ S1AHSF400W40_WLDV_2X1_882_SB
XWLDV_2X1<9> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[36] WL[37] WL[38] WL[39] 
+ S1AHSF400W40_WLDV_2X1_882_SB
XWLDV_2X1<10> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[5] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[40] WL[41] WL[42] WL[43] 
+ S1AHSF400W40_WLDV_2X1_882_SB
XWLDV_2X1<11> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[44] WL[45] WL[46] WL[47] 
+ S1AHSF400W40_WLDV_2X1_882_SB
XWLDV_2X1<12> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[6] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[48] WL[49] WL[50] WL[51] 
+ S1AHSF400W40_WLDV_2X1_882_SB
XWLDV_2X1<13> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[52] WL[53] WL[54] WL[55] 
+ S1AHSF400W40_WLDV_2X1_882_SB
XWLDV_2X1<14> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[7] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[56] WL[57] WL[58] WL[59] 
+ S1AHSF400W40_WLDV_2X1_882_SB
XWLDV_2X1<15> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[60] WL[61] WL[62] WL[63] 
+ S1AHSF400W40_WLDV_2X1_882_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_882_LD_U_64
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_882_LD_U_64 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2_SHARE 
+ PD_BUF VDDHD VDDI VSSI
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2_SHARE:B PD_BUF:B VDDHD:B 
*.PININFO VDDI:B VSSI:B
XWLDV_64X1 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI 
+ NET20[0] NET20[1] NET20[2] NET20[3] NET20[4] NET20[5] NET20[6] NET20[7] 
+ NET20[8] NET20[9] NET20[10] NET20[11] NET20[12] NET20[13] NET20[14] 
+ NET20[15] NET20[16] NET20[17] NET20[18] NET20[19] NET20[20] NET20[21] 
+ NET20[22] NET20[23] NET20[24] NET20[25] NET20[26] NET20[27] NET20[28] 
+ NET20[29] NET20[30] NET20[31] NET20[32] NET20[33] NET20[34] NET20[35] 
+ NET20[36] NET20[37] NET20[38] NET20[39] NET20[40] NET20[41] NET20[42] 
+ NET20[43] NET20[44] NET20[45] NET20[46] NET20[47] NET20[48] NET20[49] 
+ NET20[50] NET20[51] NET20[52] NET20[53] NET20[54] NET20[55] NET20[56] 
+ NET20[57] NET20[58] NET20[59] NET20[60] NET20[61] NET20[62] NET20[63] 
+ S1AHSF400W40_WLDV_64X1_882_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    WLDV_2X1_888_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_WLDV_2X1_888_SB DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1 DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[0] WL[1] WL[2] WL[3]
*.PININFO DEC_X0[0]:I DEC_X0[1]:I DEC_X0[2]:I DEC_X0[3]:I DEC_X1:I DEC_X2:I 
*.PININFO DEC_X2_SHARE:I PD_BUF:I WL[0]:O WL[1]:O WL[2]:O WL[3]:O VDDHD:B 
*.PININFO VDDI:B VSSI:B
XWLDV_0 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1 DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X2 DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[0] WL[1] S1AHSF400W40_XDRV_LA512_888_SB
XWLDV_1 DEC_X0[2] DEC_X0[3] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1 DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X2 DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[2] WL[3] S1AHSF400W40_XDRV_LA512_888_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    WLDV_64X1_888_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_WLDV_64X1_888_SB DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2 DEC_X2_SHARE PD_BUF VDDHD 
+ VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] 
+ WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] 
+ WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] 
+ WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] 
+ WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] 
+ WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63]
*.PININFO DEC_X0[0]:I DEC_X0[1]:I DEC_X0[2]:I DEC_X0[3]:I DEC_X0[4]:I 
*.PININFO DEC_X0[5]:I DEC_X0[6]:I DEC_X0[7]:I DEC_X1[0]:I DEC_X1[1]:I 
*.PININFO DEC_X1[2]:I DEC_X1[3]:I DEC_X1[4]:I DEC_X1[5]:I DEC_X1[6]:I 
*.PININFO DEC_X1[7]:I DEC_X2:I DEC_X2_SHARE:I PD_BUF:I WL[0]:O WL[1]:O WL[2]:O 
*.PININFO WL[3]:O WL[4]:O WL[5]:O WL[6]:O WL[7]:O WL[8]:O WL[9]:O WL[10]:O 
*.PININFO WL[11]:O WL[12]:O WL[13]:O WL[14]:O WL[15]:O WL[16]:O WL[17]:O 
*.PININFO WL[18]:O WL[19]:O WL[20]:O WL[21]:O WL[22]:O WL[23]:O WL[24]:O 
*.PININFO WL[25]:O WL[26]:O WL[27]:O WL[28]:O WL[29]:O WL[30]:O WL[31]:O 
*.PININFO WL[32]:O WL[33]:O WL[34]:O WL[35]:O WL[36]:O WL[37]:O WL[38]:O 
*.PININFO WL[39]:O WL[40]:O WL[41]:O WL[42]:O WL[43]:O WL[44]:O WL[45]:O 
*.PININFO WL[46]:O WL[47]:O WL[48]:O WL[49]:O WL[50]:O WL[51]:O WL[52]:O 
*.PININFO WL[53]:O WL[54]:O WL[55]:O WL[56]:O WL[57]:O WL[58]:O WL[59]:O 
*.PININFO WL[60]:O WL[61]:O WL[62]:O WL[63]:O VDDHD:B VDDI:B VSSI:B
XWLDV_2X1<0> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[0] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[0] WL[1] WL[2] WL[3] S1AHSF400W40_WLDV_2X1_888_SB
XWLDV_2X1<1> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[4] WL[5] WL[6] WL[7] S1AHSF400W40_WLDV_2X1_888_SB
XWLDV_2X1<2> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[1] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[8] WL[9] WL[10] WL[11] 
+ S1AHSF400W40_WLDV_2X1_888_SB
XWLDV_2X1<3> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[12] WL[13] WL[14] WL[15] 
+ S1AHSF400W40_WLDV_2X1_888_SB
XWLDV_2X1<4> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[2] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[16] WL[17] WL[18] WL[19] 
+ S1AHSF400W40_WLDV_2X1_888_SB
XWLDV_2X1<5> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[20] WL[21] WL[22] WL[23] 
+ S1AHSF400W40_WLDV_2X1_888_SB
XWLDV_2X1<6> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[3] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[24] WL[25] WL[26] WL[27] 
+ S1AHSF400W40_WLDV_2X1_888_SB
XWLDV_2X1<7> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[28] WL[29] WL[30] WL[31] 
+ S1AHSF400W40_WLDV_2X1_888_SB
XWLDV_2X1<8> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[4] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[32] WL[33] WL[34] WL[35] 
+ S1AHSF400W40_WLDV_2X1_888_SB
XWLDV_2X1<9> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[36] WL[37] WL[38] WL[39] 
+ S1AHSF400W40_WLDV_2X1_888_SB
XWLDV_2X1<10> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[5] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[40] WL[41] WL[42] WL[43] 
+ S1AHSF400W40_WLDV_2X1_888_SB
XWLDV_2X1<11> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[44] WL[45] WL[46] WL[47] 
+ S1AHSF400W40_WLDV_2X1_888_SB
XWLDV_2X1<12> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[6] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[48] WL[49] WL[50] WL[51] 
+ S1AHSF400W40_WLDV_2X1_888_SB
XWLDV_2X1<13> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[52] WL[53] WL[54] WL[55] 
+ S1AHSF400W40_WLDV_2X1_888_SB
XWLDV_2X1<14> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[7] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[56] WL[57] WL[58] WL[59] 
+ S1AHSF400W40_WLDV_2X1_888_SB
XWLDV_2X1<15> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[60] WL[61] WL[62] WL[63] 
+ S1AHSF400W40_WLDV_2X1_888_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_888_LD_U_384
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_888_LD_U_384 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_X2_SHARE PD_BUF VDDHD 
+ VDDI VSSI
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2[4]:B DEC_X2[5]:B DEC_X2[6]:B DEC_X2[7]:B DEC_X2_SHARE:B 
*.PININFO PD_BUF:B VDDHD:B VDDI:B VSSI:B
XWLDV_64X1 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[5] DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI 
+ NET13[0] NET13[1] NET13[2] NET13[3] NET13[4] NET13[5] NET13[6] NET13[7] 
+ NET13[8] NET13[9] NET13[10] NET13[11] NET13[12] NET13[13] NET13[14] 
+ NET13[15] NET13[16] NET13[17] NET13[18] NET13[19] NET13[20] NET13[21] 
+ NET13[22] NET13[23] NET13[24] NET13[25] NET13[26] NET13[27] NET13[28] 
+ NET13[29] NET13[30] NET13[31] NET13[32] NET13[33] NET13[34] NET13[35] 
+ NET13[36] NET13[37] NET13[38] NET13[39] NET13[40] NET13[41] NET13[42] 
+ NET13[43] NET13[44] NET13[45] NET13[46] NET13[47] NET13[48] NET13[49] 
+ NET13[50] NET13[51] NET13[52] NET13[53] NET13[54] NET13[55] NET13[56] 
+ NET13[57] NET13[58] NET13[59] NET13[60] NET13[61] NET13[62] NET13[63] 
+ S1AHSF400W40_WLDV_64X1_888_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_882_LD_U_128
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_882_LD_U_128 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2_SHARE 
+ PD_BUF VDDHD VDDI VSSI
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2_SHARE:B PD_BUF:B VDDHD:B 
*.PININFO VDDI:B VSSI:B
XWLDV_64X1 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[1] DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI 
+ NET20[0] NET20[1] NET20[2] NET20[3] NET20[4] NET20[5] NET20[6] NET20[7] 
+ NET20[8] NET20[9] NET20[10] NET20[11] NET20[12] NET20[13] NET20[14] 
+ NET20[15] NET20[16] NET20[17] NET20[18] NET20[19] NET20[20] NET20[21] 
+ NET20[22] NET20[23] NET20[24] NET20[25] NET20[26] NET20[27] NET20[28] 
+ NET20[29] NET20[30] NET20[31] NET20[32] NET20[33] NET20[34] NET20[35] 
+ NET20[36] NET20[37] NET20[38] NET20[39] NET20[40] NET20[41] NET20[42] 
+ NET20[43] NET20[44] NET20[45] NET20[46] NET20[47] NET20[48] NET20[49] 
+ NET20[50] NET20[51] NET20[52] NET20[53] NET20[54] NET20[55] NET20[56] 
+ NET20[57] NET20[58] NET20[59] NET20[60] NET20[61] NET20[62] NET20[63] 
+ S1AHSF400W40_WLDV_64X1_882_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_882_LD_U_16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_882_LD_U_16 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2_SHARE 
+ PD_BUF VDDHD VDDI VSSI
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2_SHARE:B PD_BUF:B VDDHD:B 
*.PININFO VDDI:B VSSI:B
XI39 DEC_X0[4] DEC_X0[5] NET19[0] NET19[1] NET19[2] NET19[3] NET19[4] NET19[5] 
+ DEC_X1[1] NET16[0] NET16[1] NET16[2] NET16[3] NET16[4] NET16[5] NET16[6] 
+ DEC_X2[0] NET14 DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI NET86[0] NET86[1] 
+ S1AHSF400W40_XDRV_LA512_882_SB
XI38 DEC_X0[2] DEC_X0[3] NET040[0] NET040[1] NET040[2] NET040[3] NET040[4] 
+ NET040[5] DEC_X1[1] NET28[0] NET28[1] NET28[2] NET28[3] NET28[4] NET28[5] 
+ NET28[6] DEC_X2[0] NET26 DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI NET32[0] 
+ NET32[1] S1AHSF400W40_XDRV_LA512_882_SB
XI29 DEC_X0[6] DEC_X0[7] NET43[0] NET43[1] NET43[2] NET43[3] NET43[4] NET43[5] 
+ DEC_X1[0] NET40[0] NET40[1] NET40[2] NET40[3] NET40[4] NET40[5] NET40[6] 
+ DEC_X2[0] NET38 DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI NET44[0] NET44[1] 
+ S1AHSF400W40_XDRV_LA512_882_SB
XI31 DEC_X0[4] DEC_X0[5] NET064[0] NET064[1] NET064[2] NET064[3] NET064[4] 
+ NET064[5] DEC_X1[0] NET52[0] NET52[1] NET52[2] NET52[3] NET52[4] NET52[5] 
+ NET52[6] DEC_X2[0] NET50 DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI NET56[0] 
+ NET56[1] S1AHSF400W40_XDRV_LA512_882_SB
XI34 DEC_X0[2] DEC_X0[3] NET67[0] NET67[1] NET67[2] NET67[3] NET67[4] NET67[5] 
+ DEC_X1[0] NET64[0] NET64[1] NET64[2] NET64[3] NET64[4] NET64[5] NET64[6] 
+ DEC_X2[0] NET62 DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI NET93[0] NET93[1] 
+ S1AHSF400W40_XDRV_LA512_882_SB
XI37 DEC_X0[0] DEC_X0[1] NET076[0] NET076[1] NET076[2] NET076[3] NET076[4] 
+ NET076[5] DEC_X1[1] NET76[0] NET76[1] NET76[2] NET76[3] NET76[4] NET76[5] 
+ NET76[6] DEC_X2[0] NET74 DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI NET80[0] 
+ NET80[1] S1AHSF400W40_XDRV_LA512_882_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    LD_PASS
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LD_PASS
*.PININFO
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    WLDV_2X1_884_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_WLDV_2X1_884_SB DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1 DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[0] WL[1] WL[2] WL[3]
*.PININFO DEC_X0[0]:I DEC_X0[1]:I DEC_X0[2]:I DEC_X0[3]:I DEC_X1:I DEC_X2:I 
*.PININFO DEC_X2_SHARE:I PD_BUF:I WL[0]:O WL[1]:O WL[2]:O WL[3]:O VDDHD:B 
*.PININFO VDDI:B VSSI:B
XWLDV_0 DEC_X0[0] DEC_X0[1] NET18[0] NET18[1] NET18[2] NET18[3] NET18[4] 
+ NET18[5] DEC_X1 NET20[0] NET20[1] NET20[2] NET20[3] NET20[4] NET20[5] 
+ NET20[6] DEC_X2 NET19[0] NET19[1] NET19[2] DEC_X2_SHARE PD_BUF VDDHD VDDI 
+ VSSI WL[0] WL[1] S1AHSF400W40_XDRV_LA512_884_SB
XWLDV_1 DEC_X0[2] DEC_X0[3] NET30[0] NET30[1] NET30[2] NET30[3] NET30[4] 
+ NET30[5] DEC_X1 NET32[0] NET32[1] NET32[2] NET32[3] NET32[4] NET32[5] 
+ NET32[6] DEC_X2 NET31[0] NET31[1] NET31[2] DEC_X2_SHARE PD_BUF VDDHD VDDI 
+ VSSI WL[2] WL[3] S1AHSF400W40_XDRV_LA512_884_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    WLDV_64X1_884_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_WLDV_64X1_884_SB DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2 DEC_X2_SHARE PD_BUF VDDHD 
+ VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] 
+ WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] 
+ WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] 
+ WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] 
+ WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] 
+ WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63]
*.PININFO DEC_X0[0]:I DEC_X0[1]:I DEC_X0[2]:I DEC_X0[3]:I DEC_X0[4]:I 
*.PININFO DEC_X0[5]:I DEC_X0[6]:I DEC_X0[7]:I DEC_X1[0]:I DEC_X1[1]:I 
*.PININFO DEC_X1[2]:I DEC_X1[3]:I DEC_X1[4]:I DEC_X1[5]:I DEC_X1[6]:I 
*.PININFO DEC_X1[7]:I DEC_X2:I DEC_X2_SHARE:I PD_BUF:I WL[0]:O WL[1]:O WL[2]:O 
*.PININFO WL[3]:O WL[4]:O WL[5]:O WL[6]:O WL[7]:O WL[8]:O WL[9]:O WL[10]:O 
*.PININFO WL[11]:O WL[12]:O WL[13]:O WL[14]:O WL[15]:O WL[16]:O WL[17]:O 
*.PININFO WL[18]:O WL[19]:O WL[20]:O WL[21]:O WL[22]:O WL[23]:O WL[24]:O 
*.PININFO WL[25]:O WL[26]:O WL[27]:O WL[28]:O WL[29]:O WL[30]:O WL[31]:O 
*.PININFO WL[32]:O WL[33]:O WL[34]:O WL[35]:O WL[36]:O WL[37]:O WL[38]:O 
*.PININFO WL[39]:O WL[40]:O WL[41]:O WL[42]:O WL[43]:O WL[44]:O WL[45]:O 
*.PININFO WL[46]:O WL[47]:O WL[48]:O WL[49]:O WL[50]:O WL[51]:O WL[52]:O 
*.PININFO WL[53]:O WL[54]:O WL[55]:O WL[56]:O WL[57]:O WL[58]:O WL[59]:O 
*.PININFO WL[60]:O WL[61]:O WL[62]:O WL[63]:O VDDHD:B VDDI:B VSSI:B
XWLDV_2X1<0> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[0] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[0] WL[1] WL[2] WL[3] S1AHSF400W40_WLDV_2X1_884_SB
XWLDV_2X1<1> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[4] WL[5] WL[6] WL[7] S1AHSF400W40_WLDV_2X1_884_SB
XWLDV_2X1<2> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[1] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[8] WL[9] WL[10] WL[11] 
+ S1AHSF400W40_WLDV_2X1_884_SB
XWLDV_2X1<3> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[12] WL[13] WL[14] WL[15] 
+ S1AHSF400W40_WLDV_2X1_884_SB
XWLDV_2X1<4> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[2] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[16] WL[17] WL[18] WL[19] 
+ S1AHSF400W40_WLDV_2X1_884_SB
XWLDV_2X1<5> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[20] WL[21] WL[22] WL[23] 
+ S1AHSF400W40_WLDV_2X1_884_SB
XWLDV_2X1<6> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[3] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[24] WL[25] WL[26] WL[27] 
+ S1AHSF400W40_WLDV_2X1_884_SB
XWLDV_2X1<7> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[28] WL[29] WL[30] WL[31] 
+ S1AHSF400W40_WLDV_2X1_884_SB
XWLDV_2X1<8> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[4] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[32] WL[33] WL[34] WL[35] 
+ S1AHSF400W40_WLDV_2X1_884_SB
XWLDV_2X1<9> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[36] WL[37] WL[38] WL[39] 
+ S1AHSF400W40_WLDV_2X1_884_SB
XWLDV_2X1<10> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[5] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[40] WL[41] WL[42] WL[43] 
+ S1AHSF400W40_WLDV_2X1_884_SB
XWLDV_2X1<11> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[44] WL[45] WL[46] WL[47] 
+ S1AHSF400W40_WLDV_2X1_884_SB
XWLDV_2X1<12> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[6] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[48] WL[49] WL[50] WL[51] 
+ S1AHSF400W40_WLDV_2X1_884_SB
XWLDV_2X1<13> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[52] WL[53] WL[54] WL[55] 
+ S1AHSF400W40_WLDV_2X1_884_SB
XWLDV_2X1<14> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[7] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[56] WL[57] WL[58] WL[59] 
+ S1AHSF400W40_WLDV_2X1_884_SB
XWLDV_2X1<15> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X2 
+ DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI WL[60] WL[61] WL[62] WL[63] 
+ S1AHSF400W40_WLDV_2X1_884_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_884_LD_U_256
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_884_LD_U_256 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2_SHARE:B PD_BUF:B VDDHD:B VDDI:B VSSI:B
XWLDV_64X1 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[3] DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI 
+ NET13[0] NET13[1] NET13[2] NET13[3] NET13[4] NET13[5] NET13[6] NET13[7] 
+ NET13[8] NET13[9] NET13[10] NET13[11] NET13[12] NET13[13] NET13[14] 
+ NET13[15] NET13[16] NET13[17] NET13[18] NET13[19] NET13[20] NET13[21] 
+ NET13[22] NET13[23] NET13[24] NET13[25] NET13[26] NET13[27] NET13[28] 
+ NET13[29] NET13[30] NET13[31] NET13[32] NET13[33] NET13[34] NET13[35] 
+ NET13[36] NET13[37] NET13[38] NET13[39] NET13[40] NET13[41] NET13[42] 
+ NET13[43] NET13[44] NET13[45] NET13[46] NET13[47] NET13[48] NET13[49] 
+ NET13[50] NET13[51] NET13[52] NET13[53] NET13[54] NET13[55] NET13[56] 
+ NET13[57] NET13[58] NET13[59] NET13[60] NET13[61] NET13[62] NET13[63] 
+ S1AHSF400W40_WLDV_64X1_884_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_888_LD_U_512
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_888_LD_U_512 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_X2_SHARE PD_BUF VDDHD 
+ VDDI VSSI
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2[4]:B DEC_X2[5]:B DEC_X2[6]:B DEC_X2[7]:B DEC_X2_SHARE:B 
*.PININFO PD_BUF:B VDDHD:B VDDI:B VSSI:B
XWLDV_64X1 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[7] DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI 
+ NET13[0] NET13[1] NET13[2] NET13[3] NET13[4] NET13[5] NET13[6] NET13[7] 
+ NET13[8] NET13[9] NET13[10] NET13[11] NET13[12] NET13[13] NET13[14] 
+ NET13[15] NET13[16] NET13[17] NET13[18] NET13[19] NET13[20] NET13[21] 
+ NET13[22] NET13[23] NET13[24] NET13[25] NET13[26] NET13[27] NET13[28] 
+ NET13[29] NET13[30] NET13[31] NET13[32] NET13[33] NET13[34] NET13[35] 
+ NET13[36] NET13[37] NET13[38] NET13[39] NET13[40] NET13[41] NET13[42] 
+ NET13[43] NET13[44] NET13[45] NET13[46] NET13[47] NET13[48] NET13[49] 
+ NET13[50] NET13[51] NET13[52] NET13[53] NET13[54] NET13[55] NET13[56] 
+ NET13[57] NET13[58] NET13[59] NET13[60] NET13[61] NET13[62] NET13[63] 
+ S1AHSF400W40_WLDV_64X1_888_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_BK_LD_U_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_BK_LD_U_SIM DEC_X0_BT[0] DEC_X0_BT[1] DEC_X0_BT[2] DEC_X0_BT[3] 
+ DEC_X0_BT[4] DEC_X0_BT[5] DEC_X0_BT[6] DEC_X0_BT[7] DEC_X0_TP[0] 
+ DEC_X0_TP[1] DEC_X0_TP[2] DEC_X0_TP[3] DEC_X0_TP[4] DEC_X0_TP[5] 
+ DEC_X0_TP[6] DEC_X0_TP[7] DEC_X1_BT[0] DEC_X1_BT[1] DEC_X1_BT[2] 
+ DEC_X1_BT[3] DEC_X1_BT[4] DEC_X1_BT[5] DEC_X1_BT[6] DEC_X1_BT[7] 
+ DEC_X1_TP[0] DEC_X1_TP[1] DEC_X1_TP[2] DEC_X1_TP[3] DEC_X1_TP[4] 
+ DEC_X1_TP[5] DEC_X1_TP[6] DEC_X1_TP[7] DEC_X2_BT[0] DEC_X2_BT[1] 
+ DEC_X2_BT[2] DEC_X2_BT[3] DEC_X2_BT[4] DEC_X2_BT[5] DEC_X2_BT[6] 
+ DEC_X2_BT[7] DEC_X2_SHARE_BT DEC_X2_SHARE_TP DEC_X2_TP[0] DEC_X2_TP[1] 
+ DEC_X2_TP[2] DEC_X2_TP[3] DEC_X2_TP[4] DEC_X2_TP[5] DEC_X2_TP[6] 
+ DEC_X2_TP[7] PD_BUF_BT PD_BUF_TP VDDHD VDDI VSSI
*.PININFO DEC_X0_BT[0]:B DEC_X0_BT[1]:B DEC_X0_BT[2]:B DEC_X0_BT[3]:B 
*.PININFO DEC_X0_BT[4]:B DEC_X0_BT[5]:B DEC_X0_BT[6]:B DEC_X0_BT[7]:B 
*.PININFO DEC_X0_TP[0]:B DEC_X0_TP[1]:B DEC_X0_TP[2]:B DEC_X0_TP[3]:B 
*.PININFO DEC_X0_TP[4]:B DEC_X0_TP[5]:B DEC_X0_TP[6]:B DEC_X0_TP[7]:B 
*.PININFO DEC_X1_BT[0]:B DEC_X1_BT[1]:B DEC_X1_BT[2]:B DEC_X1_BT[3]:B 
*.PININFO DEC_X1_BT[4]:B DEC_X1_BT[5]:B DEC_X1_BT[6]:B DEC_X1_BT[7]:B 
*.PININFO DEC_X1_TP[0]:B DEC_X1_TP[1]:B DEC_X1_TP[2]:B DEC_X1_TP[3]:B 
*.PININFO DEC_X1_TP[4]:B DEC_X1_TP[5]:B DEC_X1_TP[6]:B DEC_X1_TP[7]:B 
*.PININFO DEC_X2_BT[0]:B DEC_X2_BT[1]:B DEC_X2_BT[2]:B DEC_X2_BT[3]:B 
*.PININFO DEC_X2_BT[4]:B DEC_X2_BT[5]:B DEC_X2_BT[6]:B DEC_X2_BT[7]:B 
*.PININFO DEC_X2_SHARE_BT:B DEC_X2_SHARE_TP:B DEC_X2_TP[0]:B DEC_X2_TP[1]:B 
*.PININFO DEC_X2_TP[2]:B DEC_X2_TP[3]:B DEC_X2_TP[4]:B DEC_X2_TP[5]:B 
*.PININFO DEC_X2_TP[6]:B DEC_X2_TP[7]:B PD_BUF_BT:B PD_BUF_TP:B VDDHD:B VDDI:B 
*.PININFO VSSI:B
XI40 NET030[0] NET030[1] NET030[2] NET030[3] NET030[4] NET030[5] NET030[6] 
+ NET030[7] NET018[0] NET018[1] NET018[2] NET018[3] NET018[4] NET018[5] 
+ NET018[6] NET018[7] NET040[0] NET040[1] NET019 NET017 NET015 NET09 NET012 
+ S1AHSF400W40_SB_WLDV_882_LD_U_64
XI39 NET038[0] NET038[1] NET038[2] NET038[3] NET038[4] NET038[5] NET038[6] 
+ NET038[7] NET036[0] NET036[1] NET036[2] NET036[3] NET036[4] NET036[5] 
+ NET036[6] NET036[7] NET037[0] NET037[1] NET037[2] NET037[3] NET037[4] 
+ NET037[5] NET037[6] NET037[7] NET02 NET032 NET035 NET039 NET016 
+ S1AHSF400W40_SB_WLDV_888_LD_U_384
XI30 NET04[0] NET04[1] NET04[2] NET04[3] NET04[4] NET04[5] NET04[6] NET04[7] 
+ NET034[0] NET034[1] NET034[2] NET034[3] NET034[4] NET034[5] NET034[6] 
+ NET034[7] NET033[0] NET033[1] NET020 NET021 NET01 NET06 NET05 
+ S1AHSF400W40_SB_WLDV_882_LD_U_128
XI31 NET031[0] NET031[1] NET031[2] NET031[3] NET031[4] NET031[5] NET031[6] 
+ NET031[7] NET042[0] NET042[1] NET042[2] NET042[3] NET042[4] NET042[5] 
+ NET042[6] NET042[7] NET041[0] NET041[1] NET07 NET011 NET03 NET08 NET010 
+ S1AHSF400W40_SB_WLDV_882_LD_U_16
XI37  S1AHSF400W40_LD_PASS
XI34  S1AHSF400W40_LD_PASS
XI35  S1AHSF400W40_LD_PASS
XI36  S1AHSF400W40_LD_PASS
XI25 NET19[0] NET19[1] NET19[2] NET19[3] NET19[4] NET19[5] NET19[6] NET19[7] 
+ NET18[0] NET18[1] NET18[2] NET18[3] NET18[4] NET18[5] NET18[6] NET18[7] 
+ NET014[0] NET014[1] NET014[2] NET014[3] NET013 NET12 NET16 NET15 NET14 
+ S1AHSF400W40_SB_WLDV_884_LD_U_256
XI26 NET029[0] NET029[1] NET029[2] NET029[3] NET029[4] NET029[5] NET029[6] 
+ NET029[7] NET027[0] NET027[1] NET027[2] NET027[3] NET027[4] NET027[5] 
+ NET027[6] NET027[7] NET028[0] NET028[1] NET028[2] NET028[3] NET028[4] 
+ NET028[5] NET028[6] NET028[7] NET022 NET023 NET026 NET025 NET024 
+ S1AHSF400W40_SB_WLDV_888_LD_U_512
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_ARR_MCB_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_ARR_MCB_SIM BLB_BT[0] BLB_TP[0] BL_BT[0] BL_TP[0] CVDDI VDDHD VDDI 
+ VSSI WL_LT[0] WL_LT[1] WL_RT[0] WL_RT[1]
*.PININFO BLB_BT[0]:B BLB_TP[0]:B BL_BT[0]:B BL_TP[0]:B CVDDI:B VDDHD:B VDDI:B 
*.PININFO VSSI:B WL_LT[0]:B WL_LT[1]:B WL_RT[0]:B WL_RT[1]:B
XI23 NET011[0] NET011[1] NET011[2] NET011[3] NET011[4] NET011[5] NET011[6] 
+ NET011[7] NET011[8] NET011[9] NET011[10] NET011[11] NET011[12] NET011[13] 
+ NET011[14] NET011[15] NET012[0] NET012[1] NET012[2] NET012[3] NET012[4] 
+ NET012[5] NET012[6] NET012[7] NET012[8] NET012[9] NET012[10] NET012[11] 
+ NET012[12] NET012[13] NET012[14] NET012[15] NET015 NET014 NET013[0] 
+ NET013[1] S1AHSF400W40_MCB_2X16_SB_CHAR
XI22 NET017[0] NET017[1] NET017[2] NET017[3] NET017[4] NET017[5] NET017[6] 
+ NET017[7] NET016[0] NET016[1] NET016[2] NET016[3] NET016[4] NET016[5] 
+ NET016[6] NET016[7] NET020 NET019 NET018[0] NET018[1] S1AHSF400W40_MCB_2X8_SB_CHAR
XI265 NET15[0] NET15[1] NET15[2] NET15[3] NET11[0] NET11[1] NET11[2] NET11[3] 
+ NET14 NET13 NET12[0] NET12[1] S1AHSF400W40_MCB_2X4_SB_CHAR
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MCB_2X4_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_2X4_SB BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI 
+ VSSI WL[0] WL[1]
*.PININFO WL[0]:I WL[1]:I BL[0]:B BL[1]:B BL[2]:B BL[3]:B BLB[0]:B BLB[1]:B 
*.PININFO BLB[2]:B BLB[3]:B VDDI:B VSSI:B
XMCB_0<0> BL[0] BLB[0] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<1> BL[1] BLB[1] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<2> BL[2] BLB[2] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<3> BL[3] BLB[3] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_1<0> BL[0] BLB[0] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<1> BL[1] BLB[1] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<2> BL[2] BLB[2] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<3> BL[3] BLB[3] VDDI VSSI WL[1] S1AHSF400W40_MCB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    MCB_62X4_SB_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_62X4_SB_CHAR BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] 
+ VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] 
+ WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] 
+ WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] 
+ WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] 
+ WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] 
+ WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61]
*.PININFO WL[0]:I WL[1]:I WL[2]:I WL[3]:I WL[4]:I WL[5]:I WL[6]:I WL[7]:I 
*.PININFO WL[8]:I WL[9]:I WL[10]:I WL[11]:I WL[12]:I WL[13]:I WL[14]:I 
*.PININFO WL[15]:I WL[16]:I WL[17]:I WL[18]:I WL[19]:I WL[20]:I WL[21]:I 
*.PININFO WL[22]:I WL[23]:I WL[24]:I WL[25]:I WL[26]:I WL[27]:I WL[28]:I 
*.PININFO WL[29]:I WL[30]:I WL[31]:I WL[32]:I WL[33]:I WL[34]:I WL[35]:I 
*.PININFO WL[36]:I WL[37]:I WL[38]:I WL[39]:I WL[40]:I WL[41]:I WL[42]:I 
*.PININFO WL[43]:I WL[44]:I WL[45]:I WL[46]:I WL[47]:I WL[48]:I WL[49]:I 
*.PININFO WL[50]:I WL[51]:I WL[52]:I WL[53]:I WL[54]:I WL[55]:I WL[56]:I 
*.PININFO WL[57]:I WL[58]:I WL[59]:I WL[60]:I WL[61]:I BL[0]:B BL[1]:B BL[2]:B 
*.PININFO BL[3]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B VDDI:B VSSI:B
XMCB_2X4<0> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[0] WL[1] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<1> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[2] WL[3] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<2> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[4] WL[5] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<3> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[6] WL[7] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<4> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[8] WL[9] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<5> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[10] WL[11] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<6> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[12] WL[13] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<7> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[14] WL[15] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<8> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[16] WL[17] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<9> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[18] WL[19] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<10> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[20] WL[21] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<11> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[22] WL[23] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<12> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[24] WL[25] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<13> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[26] WL[27] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<14> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[28] WL[29] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<15> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[30] WL[31] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<16> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[32] WL[33] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<17> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[34] WL[35] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<18> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[36] WL[37] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<19> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[38] WL[39] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<20> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[40] WL[41] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<21> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[42] WL[43] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<22> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[44] WL[45] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<23> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[46] WL[47] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<24> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[48] WL[49] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<25> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[50] WL[51] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<26> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[52] WL[53] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<27> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[54] WL[55] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<28> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[56] WL[57] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<29> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[58] WL[59] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<30> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[60] WL[61] S1AHSF400W40_MCB_2X4_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    MCB_60X4_SB_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_60X4_SB_CHAR BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] 
+ VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] 
+ WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] 
+ WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] 
+ WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] 
+ WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] 
+ WL[55] WL[56] WL[57] WL[58] WL[59]
*.PININFO WL[0]:I WL[1]:I WL[2]:I WL[3]:I WL[4]:I WL[5]:I WL[6]:I WL[7]:I 
*.PININFO WL[8]:I WL[9]:I WL[10]:I WL[11]:I WL[12]:I WL[13]:I WL[14]:I 
*.PININFO WL[15]:I WL[16]:I WL[17]:I WL[18]:I WL[19]:I WL[20]:I WL[21]:I 
*.PININFO WL[22]:I WL[23]:I WL[24]:I WL[25]:I WL[26]:I WL[27]:I WL[28]:I 
*.PININFO WL[29]:I WL[30]:I WL[31]:I WL[32]:I WL[33]:I WL[34]:I WL[35]:I 
*.PININFO WL[36]:I WL[37]:I WL[38]:I WL[39]:I WL[40]:I WL[41]:I WL[42]:I 
*.PININFO WL[43]:I WL[44]:I WL[45]:I WL[46]:I WL[47]:I WL[48]:I WL[49]:I 
*.PININFO WL[50]:I WL[51]:I WL[52]:I WL[53]:I WL[54]:I WL[55]:I WL[56]:I 
*.PININFO WL[57]:I WL[58]:I WL[59]:I BL[0]:B BL[1]:B BL[2]:B BL[3]:B BLB[0]:B 
*.PININFO BLB[1]:B BLB[2]:B BLB[3]:B VDDI:B VSSI:B
XMCB_2X4<0> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[0] WL[1] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<1> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[2] WL[3] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<2> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[4] WL[5] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<3> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[6] WL[7] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<4> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[8] WL[9] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<5> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[10] WL[11] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<6> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[12] WL[13] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<7> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[14] WL[15] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<8> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[16] WL[17] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<9> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[18] WL[19] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<10> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[20] WL[21] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<11> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[22] WL[23] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<12> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[24] WL[25] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<13> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[26] WL[27] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<14> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[28] WL[29] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<15> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[30] WL[31] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<16> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[32] WL[33] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<17> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[34] WL[35] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<18> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[36] WL[37] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<19> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[38] WL[39] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<20> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[40] WL[41] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<21> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[42] WL[43] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<22> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[44] WL[45] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<23> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[46] WL[47] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<24> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[48] WL[49] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<25> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[50] WL[51] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<26> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[52] WL[53] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<27> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[54] WL[55] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<28> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[56] WL[57] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<29> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[58] WL[59] S1AHSF400W40_MCB_2X4_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    MCB_380X4_SB_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_380X4_SB_CHAR BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] 
+ VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] 
+ WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] 
+ WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] 
+ WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] 
+ WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] 
+ WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] WL[64] WL[65] 
+ WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] 
+ WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] 
+ WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] 
+ WL[99] WL[100] WL[101] WL[102] WL[103] WL[104] WL[105] WL[106] WL[107] 
+ WL[108] WL[109] WL[110] WL[111] WL[112] WL[113] WL[114] WL[115] WL[116] 
+ WL[117] WL[118] WL[119] WL[120] WL[121] WL[122] WL[123] WL[124] WL[125] 
+ WL[126] WL[127] WL[128] WL[129] WL[130] WL[131] WL[132] WL[133] WL[134] 
+ WL[135] WL[136] WL[137] WL[138] WL[139] WL[140] WL[141] WL[142] WL[143] 
+ WL[144] WL[145] WL[146] WL[147] WL[148] WL[149] WL[150] WL[151] WL[152] 
+ WL[153] WL[154] WL[155] WL[156] WL[157] WL[158] WL[159] WL[160] WL[161] 
+ WL[162] WL[163] WL[164] WL[165] WL[166] WL[167] WL[168] WL[169] WL[170] 
+ WL[171] WL[172] WL[173] WL[174] WL[175] WL[176] WL[177] WL[178] WL[179] 
+ WL[180] WL[181] WL[182] WL[183] WL[184] WL[185] WL[186] WL[187] WL[188] 
+ WL[189] WL[190] WL[191] WL[192] WL[193] WL[194] WL[195] WL[196] WL[197] 
+ WL[198] WL[199] WL[200] WL[201] WL[202] WL[203] WL[204] WL[205] WL[206] 
+ WL[207] WL[208] WL[209] WL[210] WL[211] WL[212] WL[213] WL[214] WL[215] 
+ WL[216] WL[217] WL[218] WL[219] WL[220] WL[221] WL[222] WL[223] WL[224] 
+ WL[225] WL[226] WL[227] WL[228] WL[229] WL[230] WL[231] WL[232] WL[233] 
+ WL[234] WL[235] WL[236] WL[237] WL[238] WL[239] WL[240] WL[241] WL[242] 
+ WL[243] WL[244] WL[245] WL[246] WL[247] WL[248] WL[249] WL[250] WL[251] 
+ WL[252] WL[253] WL[254] WL[255] WL[256] WL[257] WL[258] WL[259] WL[260] 
+ WL[261] WL[262] WL[263] WL[264] WL[265] WL[266] WL[267] WL[268] WL[269] 
+ WL[270] WL[271] WL[272] WL[273] WL[274] WL[275] WL[276] WL[277] WL[278] 
+ WL[279] WL[280] WL[281] WL[282] WL[283] WL[284] WL[285] WL[286] WL[287] 
+ WL[288] WL[289] WL[290] WL[291] WL[292] WL[293] WL[294] WL[295] WL[296] 
+ WL[297] WL[298] WL[299] WL[300] WL[301] WL[302] WL[303] WL[304] WL[305] 
+ WL[306] WL[307] WL[308] WL[309] WL[310] WL[311] WL[312] WL[313] WL[314] 
+ WL[315] WL[316] WL[317] WL[318] WL[319] WL[320] WL[321] WL[322] WL[323] 
+ WL[324] WL[325] WL[326] WL[327] WL[328] WL[329] WL[330] WL[331] WL[332] 
+ WL[333] WL[334] WL[335] WL[336] WL[337] WL[338] WL[339] WL[340] WL[341] 
+ WL[342] WL[343] WL[344] WL[345] WL[346] WL[347] WL[348] WL[349] WL[350] 
+ WL[351] WL[352] WL[353] WL[354] WL[355] WL[356] WL[357] WL[358] WL[359] 
+ WL[360] WL[361] WL[362] WL[363] WL[364] WL[365] WL[366] WL[367] WL[368] 
+ WL[369] WL[370] WL[371] WL[372] WL[373] WL[374] WL[375] WL[376] WL[377] 
+ WL[378] WL[379]
*.PININFO WL[0]:I WL[1]:I WL[2]:I WL[3]:I WL[4]:I WL[5]:I WL[6]:I WL[7]:I 
*.PININFO WL[8]:I WL[9]:I WL[10]:I WL[11]:I WL[12]:I WL[13]:I WL[14]:I 
*.PININFO WL[15]:I WL[16]:I WL[17]:I WL[18]:I WL[19]:I WL[20]:I WL[21]:I 
*.PININFO WL[22]:I WL[23]:I WL[24]:I WL[25]:I WL[26]:I WL[27]:I WL[28]:I 
*.PININFO WL[29]:I WL[30]:I WL[31]:I WL[32]:I WL[33]:I WL[34]:I WL[35]:I 
*.PININFO WL[36]:I WL[37]:I WL[38]:I WL[39]:I WL[40]:I WL[41]:I WL[42]:I 
*.PININFO WL[43]:I WL[44]:I WL[45]:I WL[46]:I WL[47]:I WL[48]:I WL[49]:I 
*.PININFO WL[50]:I WL[51]:I WL[52]:I WL[53]:I WL[54]:I WL[55]:I WL[56]:I 
*.PININFO WL[57]:I WL[58]:I WL[59]:I WL[60]:I WL[61]:I WL[62]:I WL[63]:I 
*.PININFO WL[64]:I WL[65]:I WL[66]:I WL[67]:I WL[68]:I WL[69]:I WL[70]:I 
*.PININFO WL[71]:I WL[72]:I WL[73]:I WL[74]:I WL[75]:I WL[76]:I WL[77]:I 
*.PININFO WL[78]:I WL[79]:I WL[80]:I WL[81]:I WL[82]:I WL[83]:I WL[84]:I 
*.PININFO WL[85]:I WL[86]:I WL[87]:I WL[88]:I WL[89]:I WL[90]:I WL[91]:I 
*.PININFO WL[92]:I WL[93]:I WL[94]:I WL[95]:I WL[96]:I WL[97]:I WL[98]:I 
*.PININFO WL[99]:I WL[100]:I WL[101]:I WL[102]:I WL[103]:I WL[104]:I WL[105]:I 
*.PININFO WL[106]:I WL[107]:I WL[108]:I WL[109]:I WL[110]:I WL[111]:I 
*.PININFO WL[112]:I WL[113]:I WL[114]:I WL[115]:I WL[116]:I WL[117]:I 
*.PININFO WL[118]:I WL[119]:I WL[120]:I WL[121]:I WL[122]:I WL[123]:I 
*.PININFO WL[124]:I WL[125]:I WL[126]:I WL[127]:I WL[128]:I WL[129]:I 
*.PININFO WL[130]:I WL[131]:I WL[132]:I WL[133]:I WL[134]:I WL[135]:I 
*.PININFO WL[136]:I WL[137]:I WL[138]:I WL[139]:I WL[140]:I WL[141]:I 
*.PININFO WL[142]:I WL[143]:I WL[144]:I WL[145]:I WL[146]:I WL[147]:I 
*.PININFO WL[148]:I WL[149]:I WL[150]:I WL[151]:I WL[152]:I WL[153]:I 
*.PININFO WL[154]:I WL[155]:I WL[156]:I WL[157]:I WL[158]:I WL[159]:I 
*.PININFO WL[160]:I WL[161]:I WL[162]:I WL[163]:I WL[164]:I WL[165]:I 
*.PININFO WL[166]:I WL[167]:I WL[168]:I WL[169]:I WL[170]:I WL[171]:I 
*.PININFO WL[172]:I WL[173]:I WL[174]:I WL[175]:I WL[176]:I WL[177]:I 
*.PININFO WL[178]:I WL[179]:I WL[180]:I WL[181]:I WL[182]:I WL[183]:I 
*.PININFO WL[184]:I WL[185]:I WL[186]:I WL[187]:I WL[188]:I WL[189]:I 
*.PININFO WL[190]:I WL[191]:I WL[192]:I WL[193]:I WL[194]:I WL[195]:I 
*.PININFO WL[196]:I WL[197]:I WL[198]:I WL[199]:I WL[200]:I WL[201]:I 
*.PININFO WL[202]:I WL[203]:I WL[204]:I WL[205]:I WL[206]:I WL[207]:I 
*.PININFO WL[208]:I WL[209]:I WL[210]:I WL[211]:I WL[212]:I WL[213]:I 
*.PININFO WL[214]:I WL[215]:I WL[216]:I WL[217]:I WL[218]:I WL[219]:I 
*.PININFO WL[220]:I WL[221]:I WL[222]:I WL[223]:I WL[224]:I WL[225]:I 
*.PININFO WL[226]:I WL[227]:I WL[228]:I WL[229]:I WL[230]:I WL[231]:I 
*.PININFO WL[232]:I WL[233]:I WL[234]:I WL[235]:I WL[236]:I WL[237]:I 
*.PININFO WL[238]:I WL[239]:I WL[240]:I WL[241]:I WL[242]:I WL[243]:I 
*.PININFO WL[244]:I WL[245]:I WL[246]:I WL[247]:I WL[248]:I WL[249]:I 
*.PININFO WL[250]:I WL[251]:I WL[252]:I WL[253]:I WL[254]:I WL[255]:I 
*.PININFO WL[256]:I WL[257]:I WL[258]:I WL[259]:I WL[260]:I WL[261]:I 
*.PININFO WL[262]:I WL[263]:I WL[264]:I WL[265]:I WL[266]:I WL[267]:I 
*.PININFO WL[268]:I WL[269]:I WL[270]:I WL[271]:I WL[272]:I WL[273]:I 
*.PININFO WL[274]:I WL[275]:I WL[276]:I WL[277]:I WL[278]:I WL[279]:I 
*.PININFO WL[280]:I WL[281]:I WL[282]:I WL[283]:I WL[284]:I WL[285]:I 
*.PININFO WL[286]:I WL[287]:I WL[288]:I WL[289]:I WL[290]:I WL[291]:I 
*.PININFO WL[292]:I WL[293]:I WL[294]:I WL[295]:I WL[296]:I WL[297]:I 
*.PININFO WL[298]:I WL[299]:I WL[300]:I WL[301]:I WL[302]:I WL[303]:I 
*.PININFO WL[304]:I WL[305]:I WL[306]:I WL[307]:I WL[308]:I WL[309]:I 
*.PININFO WL[310]:I WL[311]:I WL[312]:I WL[313]:I WL[314]:I WL[315]:I 
*.PININFO WL[316]:I WL[317]:I WL[318]:I WL[319]:I WL[320]:I WL[321]:I 
*.PININFO WL[322]:I WL[323]:I WL[324]:I WL[325]:I WL[326]:I WL[327]:I 
*.PININFO WL[328]:I WL[329]:I WL[330]:I WL[331]:I WL[332]:I WL[333]:I 
*.PININFO WL[334]:I WL[335]:I WL[336]:I WL[337]:I WL[338]:I WL[339]:I 
*.PININFO WL[340]:I WL[341]:I WL[342]:I WL[343]:I WL[344]:I WL[345]:I 
*.PININFO WL[346]:I WL[347]:I WL[348]:I WL[349]:I WL[350]:I WL[351]:I 
*.PININFO WL[352]:I WL[353]:I WL[354]:I WL[355]:I WL[356]:I WL[357]:I 
*.PININFO WL[358]:I WL[359]:I WL[360]:I WL[361]:I WL[362]:I WL[363]:I 
*.PININFO WL[364]:I WL[365]:I WL[366]:I WL[367]:I WL[368]:I WL[369]:I 
*.PININFO WL[370]:I WL[371]:I WL[372]:I WL[373]:I WL[374]:I WL[375]:I 
*.PININFO WL[376]:I WL[377]:I WL[378]:I WL[379]:I BL[0]:B BL[1]:B BL[2]:B 
*.PININFO BL[3]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B VDDI:B VSSI:B
XMCB_2X4<0> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[0] WL[1] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<1> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[2] WL[3] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<2> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[4] WL[5] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<3> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[6] WL[7] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<4> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[8] WL[9] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<5> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[10] WL[11] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<6> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[12] WL[13] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<7> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[14] WL[15] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<8> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[16] WL[17] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<9> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[18] WL[19] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<10> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[20] WL[21] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<11> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[22] WL[23] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<12> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[24] WL[25] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<13> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[26] WL[27] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<14> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[28] WL[29] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<15> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[30] WL[31] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<16> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[32] WL[33] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<17> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[34] WL[35] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<18> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[36] WL[37] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<19> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[38] WL[39] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<20> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[40] WL[41] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<21> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[42] WL[43] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<22> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[44] WL[45] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<23> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[46] WL[47] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<24> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[48] WL[49] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<25> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[50] WL[51] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<26> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[52] WL[53] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<27> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[54] WL[55] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<28> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[56] WL[57] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<29> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[58] WL[59] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<30> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[60] WL[61] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<31> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[62] WL[63] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<32> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[64] WL[65] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<33> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[66] WL[67] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<34> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[68] WL[69] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<35> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[70] WL[71] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<36> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[72] WL[73] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<37> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[74] WL[75] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<38> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[76] WL[77] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<39> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[78] WL[79] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<40> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[80] WL[81] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<41> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[82] WL[83] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<42> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[84] WL[85] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<43> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[86] WL[87] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<44> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[88] WL[89] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<45> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[90] WL[91] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<46> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[92] WL[93] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<47> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[94] WL[95] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<48> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[96] WL[97] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<49> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[98] WL[99] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<50> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[100] WL[101] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<51> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[102] WL[103] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<52> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[104] WL[105] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<53> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[106] WL[107] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<54> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[108] WL[109] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<55> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[110] WL[111] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<56> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[112] WL[113] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<57> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[114] WL[115] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<58> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[116] WL[117] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<59> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[118] WL[119] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<60> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[120] WL[121] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<61> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[122] WL[123] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<62> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[124] WL[125] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<63> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[126] WL[127] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<64> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[128] WL[129] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<65> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[130] WL[131] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<66> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[132] WL[133] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<67> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[134] WL[135] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<68> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[136] WL[137] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<69> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[138] WL[139] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<70> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[140] WL[141] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<71> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[142] WL[143] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<72> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[144] WL[145] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<73> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[146] WL[147] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<74> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[148] WL[149] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<75> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[150] WL[151] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<76> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[152] WL[153] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<77> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[154] WL[155] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<78> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[156] WL[157] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<79> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[158] WL[159] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<80> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[160] WL[161] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<81> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[162] WL[163] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<82> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[164] WL[165] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<83> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[166] WL[167] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<84> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[168] WL[169] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<85> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[170] WL[171] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<86> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[172] WL[173] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<87> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[174] WL[175] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<88> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[176] WL[177] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<89> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[178] WL[179] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<90> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[180] WL[181] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<91> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[182] WL[183] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<92> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[184] WL[185] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<93> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[186] WL[187] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<94> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[188] WL[189] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<95> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[190] WL[191] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<96> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[192] WL[193] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<97> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[194] WL[195] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<98> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[196] WL[197] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<99> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[198] WL[199] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<100> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[200] WL[201] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<101> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[202] WL[203] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<102> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[204] WL[205] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<103> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[206] WL[207] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<104> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[208] WL[209] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<105> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[210] WL[211] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<106> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[212] WL[213] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<107> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[214] WL[215] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<108> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[216] WL[217] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<109> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[218] WL[219] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<110> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[220] WL[221] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<111> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[222] WL[223] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<112> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[224] WL[225] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<113> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[226] WL[227] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<114> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[228] WL[229] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<115> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[230] WL[231] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<116> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[232] WL[233] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<117> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[234] WL[235] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<118> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[236] WL[237] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<119> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[238] WL[239] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<120> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[240] WL[241] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<121> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[242] WL[243] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<122> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[244] WL[245] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<123> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[246] WL[247] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<124> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[248] WL[249] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<125> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[250] WL[251] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<126> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[252] WL[253] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<127> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[254] WL[255] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<128> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[256] WL[257] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<129> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[258] WL[259] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<130> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[260] WL[261] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<131> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[262] WL[263] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<132> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[264] WL[265] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<133> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[266] WL[267] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<134> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[268] WL[269] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<135> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[270] WL[271] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<136> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[272] WL[273] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<137> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[274] WL[275] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<138> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[276] WL[277] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<139> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[278] WL[279] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<140> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[280] WL[281] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<141> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[282] WL[283] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<142> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[284] WL[285] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<143> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[286] WL[287] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<144> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[288] WL[289] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<145> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[290] WL[291] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<146> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[292] WL[293] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<147> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[294] WL[295] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<148> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[296] WL[297] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<149> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[298] WL[299] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<150> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[300] WL[301] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<151> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[302] WL[303] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<152> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[304] WL[305] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<153> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[306] WL[307] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<154> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[308] WL[309] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<155> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[310] WL[311] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<156> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[312] WL[313] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<157> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[314] WL[315] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<158> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[316] WL[317] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<159> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[318] WL[319] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<160> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[320] WL[321] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<161> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[322] WL[323] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<162> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[324] WL[325] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<163> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[326] WL[327] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<164> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[328] WL[329] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<165> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[330] WL[331] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<166> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[332] WL[333] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<167> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[334] WL[335] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<168> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[336] WL[337] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<169> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[338] WL[339] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<170> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[340] WL[341] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<171> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[342] WL[343] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<172> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[344] WL[345] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<173> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[346] WL[347] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<174> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[348] WL[349] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<175> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[350] WL[351] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<176> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[352] WL[353] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<177> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[354] WL[355] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<178> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[356] WL[357] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<179> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[358] WL[359] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<180> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[360] WL[361] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<181> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[362] WL[363] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<182> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[364] WL[365] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<183> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[366] WL[367] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<184> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[368] WL[369] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<185> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[370] WL[371] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<186> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[372] WL[373] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<187> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[374] WL[375] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<188> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[376] WL[377] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<189> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[378] WL[379] S1AHSF400W40_MCB_2X4_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    MCB_382X4_SB_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_382X4_SB_CHAR BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] 
+ VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] 
+ WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] 
+ WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] 
+ WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] 
+ WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] 
+ WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] WL[64] WL[65] 
+ WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] 
+ WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] 
+ WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] 
+ WL[99] WL[100] WL[101] WL[102] WL[103] WL[104] WL[105] WL[106] WL[107] 
+ WL[108] WL[109] WL[110] WL[111] WL[112] WL[113] WL[114] WL[115] WL[116] 
+ WL[117] WL[118] WL[119] WL[120] WL[121] WL[122] WL[123] WL[124] WL[125] 
+ WL[126] WL[127] WL[128] WL[129] WL[130] WL[131] WL[132] WL[133] WL[134] 
+ WL[135] WL[136] WL[137] WL[138] WL[139] WL[140] WL[141] WL[142] WL[143] 
+ WL[144] WL[145] WL[146] WL[147] WL[148] WL[149] WL[150] WL[151] WL[152] 
+ WL[153] WL[154] WL[155] WL[156] WL[157] WL[158] WL[159] WL[160] WL[161] 
+ WL[162] WL[163] WL[164] WL[165] WL[166] WL[167] WL[168] WL[169] WL[170] 
+ WL[171] WL[172] WL[173] WL[174] WL[175] WL[176] WL[177] WL[178] WL[179] 
+ WL[180] WL[181] WL[182] WL[183] WL[184] WL[185] WL[186] WL[187] WL[188] 
+ WL[189] WL[190] WL[191] WL[192] WL[193] WL[194] WL[195] WL[196] WL[197] 
+ WL[198] WL[199] WL[200] WL[201] WL[202] WL[203] WL[204] WL[205] WL[206] 
+ WL[207] WL[208] WL[209] WL[210] WL[211] WL[212] WL[213] WL[214] WL[215] 
+ WL[216] WL[217] WL[218] WL[219] WL[220] WL[221] WL[222] WL[223] WL[224] 
+ WL[225] WL[226] WL[227] WL[228] WL[229] WL[230] WL[231] WL[232] WL[233] 
+ WL[234] WL[235] WL[236] WL[237] WL[238] WL[239] WL[240] WL[241] WL[242] 
+ WL[243] WL[244] WL[245] WL[246] WL[247] WL[248] WL[249] WL[250] WL[251] 
+ WL[252] WL[253] WL[254] WL[255] WL[256] WL[257] WL[258] WL[259] WL[260] 
+ WL[261] WL[262] WL[263] WL[264] WL[265] WL[266] WL[267] WL[268] WL[269] 
+ WL[270] WL[271] WL[272] WL[273] WL[274] WL[275] WL[276] WL[277] WL[278] 
+ WL[279] WL[280] WL[281] WL[282] WL[283] WL[284] WL[285] WL[286] WL[287] 
+ WL[288] WL[289] WL[290] WL[291] WL[292] WL[293] WL[294] WL[295] WL[296] 
+ WL[297] WL[298] WL[299] WL[300] WL[301] WL[302] WL[303] WL[304] WL[305] 
+ WL[306] WL[307] WL[308] WL[309] WL[310] WL[311] WL[312] WL[313] WL[314] 
+ WL[315] WL[316] WL[317] WL[318] WL[319] WL[320] WL[321] WL[322] WL[323] 
+ WL[324] WL[325] WL[326] WL[327] WL[328] WL[329] WL[330] WL[331] WL[332] 
+ WL[333] WL[334] WL[335] WL[336] WL[337] WL[338] WL[339] WL[340] WL[341] 
+ WL[342] WL[343] WL[344] WL[345] WL[346] WL[347] WL[348] WL[349] WL[350] 
+ WL[351] WL[352] WL[353] WL[354] WL[355] WL[356] WL[357] WL[358] WL[359] 
+ WL[360] WL[361] WL[362] WL[363] WL[364] WL[365] WL[366] WL[367] WL[368] 
+ WL[369] WL[370] WL[371] WL[372] WL[373] WL[374] WL[375] WL[376] WL[377] 
+ WL[378] WL[379] WL[380] WL[381]
*.PININFO WL[0]:I WL[1]:I WL[2]:I WL[3]:I WL[4]:I WL[5]:I WL[6]:I WL[7]:I 
*.PININFO WL[8]:I WL[9]:I WL[10]:I WL[11]:I WL[12]:I WL[13]:I WL[14]:I 
*.PININFO WL[15]:I WL[16]:I WL[17]:I WL[18]:I WL[19]:I WL[20]:I WL[21]:I 
*.PININFO WL[22]:I WL[23]:I WL[24]:I WL[25]:I WL[26]:I WL[27]:I WL[28]:I 
*.PININFO WL[29]:I WL[30]:I WL[31]:I WL[32]:I WL[33]:I WL[34]:I WL[35]:I 
*.PININFO WL[36]:I WL[37]:I WL[38]:I WL[39]:I WL[40]:I WL[41]:I WL[42]:I 
*.PININFO WL[43]:I WL[44]:I WL[45]:I WL[46]:I WL[47]:I WL[48]:I WL[49]:I 
*.PININFO WL[50]:I WL[51]:I WL[52]:I WL[53]:I WL[54]:I WL[55]:I WL[56]:I 
*.PININFO WL[57]:I WL[58]:I WL[59]:I WL[60]:I WL[61]:I WL[62]:I WL[63]:I 
*.PININFO WL[64]:I WL[65]:I WL[66]:I WL[67]:I WL[68]:I WL[69]:I WL[70]:I 
*.PININFO WL[71]:I WL[72]:I WL[73]:I WL[74]:I WL[75]:I WL[76]:I WL[77]:I 
*.PININFO WL[78]:I WL[79]:I WL[80]:I WL[81]:I WL[82]:I WL[83]:I WL[84]:I 
*.PININFO WL[85]:I WL[86]:I WL[87]:I WL[88]:I WL[89]:I WL[90]:I WL[91]:I 
*.PININFO WL[92]:I WL[93]:I WL[94]:I WL[95]:I WL[96]:I WL[97]:I WL[98]:I 
*.PININFO WL[99]:I WL[100]:I WL[101]:I WL[102]:I WL[103]:I WL[104]:I WL[105]:I 
*.PININFO WL[106]:I WL[107]:I WL[108]:I WL[109]:I WL[110]:I WL[111]:I 
*.PININFO WL[112]:I WL[113]:I WL[114]:I WL[115]:I WL[116]:I WL[117]:I 
*.PININFO WL[118]:I WL[119]:I WL[120]:I WL[121]:I WL[122]:I WL[123]:I 
*.PININFO WL[124]:I WL[125]:I WL[126]:I WL[127]:I WL[128]:I WL[129]:I 
*.PININFO WL[130]:I WL[131]:I WL[132]:I WL[133]:I WL[134]:I WL[135]:I 
*.PININFO WL[136]:I WL[137]:I WL[138]:I WL[139]:I WL[140]:I WL[141]:I 
*.PININFO WL[142]:I WL[143]:I WL[144]:I WL[145]:I WL[146]:I WL[147]:I 
*.PININFO WL[148]:I WL[149]:I WL[150]:I WL[151]:I WL[152]:I WL[153]:I 
*.PININFO WL[154]:I WL[155]:I WL[156]:I WL[157]:I WL[158]:I WL[159]:I 
*.PININFO WL[160]:I WL[161]:I WL[162]:I WL[163]:I WL[164]:I WL[165]:I 
*.PININFO WL[166]:I WL[167]:I WL[168]:I WL[169]:I WL[170]:I WL[171]:I 
*.PININFO WL[172]:I WL[173]:I WL[174]:I WL[175]:I WL[176]:I WL[177]:I 
*.PININFO WL[178]:I WL[179]:I WL[180]:I WL[181]:I WL[182]:I WL[183]:I 
*.PININFO WL[184]:I WL[185]:I WL[186]:I WL[187]:I WL[188]:I WL[189]:I 
*.PININFO WL[190]:I WL[191]:I WL[192]:I WL[193]:I WL[194]:I WL[195]:I 
*.PININFO WL[196]:I WL[197]:I WL[198]:I WL[199]:I WL[200]:I WL[201]:I 
*.PININFO WL[202]:I WL[203]:I WL[204]:I WL[205]:I WL[206]:I WL[207]:I 
*.PININFO WL[208]:I WL[209]:I WL[210]:I WL[211]:I WL[212]:I WL[213]:I 
*.PININFO WL[214]:I WL[215]:I WL[216]:I WL[217]:I WL[218]:I WL[219]:I 
*.PININFO WL[220]:I WL[221]:I WL[222]:I WL[223]:I WL[224]:I WL[225]:I 
*.PININFO WL[226]:I WL[227]:I WL[228]:I WL[229]:I WL[230]:I WL[231]:I 
*.PININFO WL[232]:I WL[233]:I WL[234]:I WL[235]:I WL[236]:I WL[237]:I 
*.PININFO WL[238]:I WL[239]:I WL[240]:I WL[241]:I WL[242]:I WL[243]:I 
*.PININFO WL[244]:I WL[245]:I WL[246]:I WL[247]:I WL[248]:I WL[249]:I 
*.PININFO WL[250]:I WL[251]:I WL[252]:I WL[253]:I WL[254]:I WL[255]:I 
*.PININFO WL[256]:I WL[257]:I WL[258]:I WL[259]:I WL[260]:I WL[261]:I 
*.PININFO WL[262]:I WL[263]:I WL[264]:I WL[265]:I WL[266]:I WL[267]:I 
*.PININFO WL[268]:I WL[269]:I WL[270]:I WL[271]:I WL[272]:I WL[273]:I 
*.PININFO WL[274]:I WL[275]:I WL[276]:I WL[277]:I WL[278]:I WL[279]:I 
*.PININFO WL[280]:I WL[281]:I WL[282]:I WL[283]:I WL[284]:I WL[285]:I 
*.PININFO WL[286]:I WL[287]:I WL[288]:I WL[289]:I WL[290]:I WL[291]:I 
*.PININFO WL[292]:I WL[293]:I WL[294]:I WL[295]:I WL[296]:I WL[297]:I 
*.PININFO WL[298]:I WL[299]:I WL[300]:I WL[301]:I WL[302]:I WL[303]:I 
*.PININFO WL[304]:I WL[305]:I WL[306]:I WL[307]:I WL[308]:I WL[309]:I 
*.PININFO WL[310]:I WL[311]:I WL[312]:I WL[313]:I WL[314]:I WL[315]:I 
*.PININFO WL[316]:I WL[317]:I WL[318]:I WL[319]:I WL[320]:I WL[321]:I 
*.PININFO WL[322]:I WL[323]:I WL[324]:I WL[325]:I WL[326]:I WL[327]:I 
*.PININFO WL[328]:I WL[329]:I WL[330]:I WL[331]:I WL[332]:I WL[333]:I 
*.PININFO WL[334]:I WL[335]:I WL[336]:I WL[337]:I WL[338]:I WL[339]:I 
*.PININFO WL[340]:I WL[341]:I WL[342]:I WL[343]:I WL[344]:I WL[345]:I 
*.PININFO WL[346]:I WL[347]:I WL[348]:I WL[349]:I WL[350]:I WL[351]:I 
*.PININFO WL[352]:I WL[353]:I WL[354]:I WL[355]:I WL[356]:I WL[357]:I 
*.PININFO WL[358]:I WL[359]:I WL[360]:I WL[361]:I WL[362]:I WL[363]:I 
*.PININFO WL[364]:I WL[365]:I WL[366]:I WL[367]:I WL[368]:I WL[369]:I 
*.PININFO WL[370]:I WL[371]:I WL[372]:I WL[373]:I WL[374]:I WL[375]:I 
*.PININFO WL[376]:I WL[377]:I WL[378]:I WL[379]:I WL[380]:I WL[381]:I BL[0]:B 
*.PININFO BL[1]:B BL[2]:B BL[3]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B VDDI:B 
*.PININFO VSSI:B
XMCB_2X4<0> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[0] WL[1] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<1> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[2] WL[3] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<2> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[4] WL[5] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<3> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[6] WL[7] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<4> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[8] WL[9] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<5> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[10] WL[11] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<6> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[12] WL[13] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<7> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[14] WL[15] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<8> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[16] WL[17] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<9> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[18] WL[19] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<10> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[20] WL[21] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<11> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[22] WL[23] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<12> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[24] WL[25] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<13> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[26] WL[27] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<14> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[28] WL[29] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<15> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[30] WL[31] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<16> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[32] WL[33] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<17> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[34] WL[35] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<18> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[36] WL[37] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<19> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[38] WL[39] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<20> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[40] WL[41] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<21> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[42] WL[43] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<22> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[44] WL[45] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<23> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[46] WL[47] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<24> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[48] WL[49] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<25> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[50] WL[51] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<26> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[52] WL[53] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<27> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[54] WL[55] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<28> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[56] WL[57] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<29> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[58] WL[59] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<30> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[60] WL[61] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<31> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[62] WL[63] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<32> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[64] WL[65] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<33> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[66] WL[67] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<34> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[68] WL[69] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<35> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[70] WL[71] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<36> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[72] WL[73] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<37> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[74] WL[75] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<38> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[76] WL[77] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<39> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[78] WL[79] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<40> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[80] WL[81] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<41> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[82] WL[83] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<42> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[84] WL[85] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<43> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[86] WL[87] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<44> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[88] WL[89] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<45> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[90] WL[91] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<46> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[92] WL[93] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<47> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[94] WL[95] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<48> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[96] WL[97] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<49> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[98] WL[99] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<50> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[100] WL[101] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<51> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[102] WL[103] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<52> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[104] WL[105] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<53> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[106] WL[107] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<54> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[108] WL[109] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<55> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[110] WL[111] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<56> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[112] WL[113] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<57> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[114] WL[115] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<58> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[116] WL[117] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<59> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[118] WL[119] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<60> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[120] WL[121] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<61> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[122] WL[123] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<62> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[124] WL[125] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<63> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[126] WL[127] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<64> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[128] WL[129] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<65> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[130] WL[131] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<66> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[132] WL[133] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<67> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[134] WL[135] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<68> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[136] WL[137] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<69> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[138] WL[139] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<70> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[140] WL[141] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<71> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[142] WL[143] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<72> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[144] WL[145] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<73> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[146] WL[147] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<74> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[148] WL[149] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<75> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[150] WL[151] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<76> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[152] WL[153] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<77> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[154] WL[155] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<78> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[156] WL[157] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<79> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[158] WL[159] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<80> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[160] WL[161] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<81> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[162] WL[163] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<82> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[164] WL[165] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<83> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[166] WL[167] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<84> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[168] WL[169] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<85> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[170] WL[171] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<86> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[172] WL[173] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<87> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[174] WL[175] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<88> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[176] WL[177] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<89> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[178] WL[179] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<90> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[180] WL[181] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<91> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[182] WL[183] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<92> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[184] WL[185] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<93> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[186] WL[187] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<94> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[188] WL[189] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<95> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[190] WL[191] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<96> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[192] WL[193] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<97> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[194] WL[195] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<98> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[196] WL[197] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<99> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[198] WL[199] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<100> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[200] WL[201] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<101> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[202] WL[203] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<102> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[204] WL[205] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<103> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[206] WL[207] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<104> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[208] WL[209] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<105> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[210] WL[211] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<106> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[212] WL[213] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<107> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[214] WL[215] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<108> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[216] WL[217] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<109> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[218] WL[219] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<110> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[220] WL[221] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<111> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[222] WL[223] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<112> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[224] WL[225] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<113> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[226] WL[227] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<114> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[228] WL[229] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<115> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[230] WL[231] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<116> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[232] WL[233] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<117> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[234] WL[235] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<118> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[236] WL[237] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<119> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[238] WL[239] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<120> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[240] WL[241] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<121> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[242] WL[243] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<122> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[244] WL[245] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<123> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[246] WL[247] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<124> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[248] WL[249] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<125> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[250] WL[251] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<126> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[252] WL[253] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<127> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[254] WL[255] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<128> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[256] WL[257] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<129> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[258] WL[259] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<130> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[260] WL[261] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<131> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[262] WL[263] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<132> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[264] WL[265] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<133> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[266] WL[267] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<134> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[268] WL[269] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<135> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[270] WL[271] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<136> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[272] WL[273] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<137> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[274] WL[275] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<138> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[276] WL[277] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<139> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[278] WL[279] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<140> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[280] WL[281] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<141> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[282] WL[283] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<142> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[284] WL[285] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<143> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[286] WL[287] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<144> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[288] WL[289] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<145> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[290] WL[291] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<146> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[292] WL[293] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<147> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[294] WL[295] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<148> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[296] WL[297] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<149> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[298] WL[299] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<150> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[300] WL[301] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<151> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[302] WL[303] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<152> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[304] WL[305] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<153> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[306] WL[307] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<154> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[308] WL[309] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<155> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[310] WL[311] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<156> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[312] WL[313] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<157> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[314] WL[315] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<158> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[316] WL[317] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<159> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[318] WL[319] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<160> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[320] WL[321] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<161> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[322] WL[323] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<162> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[324] WL[325] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<163> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[326] WL[327] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<164> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[328] WL[329] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<165> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[330] WL[331] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<166> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[332] WL[333] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<167> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[334] WL[335] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<168> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[336] WL[337] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<169> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[338] WL[339] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<170> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[340] WL[341] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<171> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[342] WL[343] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<172> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[344] WL[345] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<173> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[346] WL[347] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<174> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[348] WL[349] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<175> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[350] WL[351] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<176> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[352] WL[353] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<177> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[354] WL[355] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<178> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[356] WL[357] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<179> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[358] WL[359] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<180> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[360] WL[361] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<181> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[362] WL[363] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<182> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[364] WL[365] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<183> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[366] WL[367] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<184> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[368] WL[369] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<185> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[370] WL[371] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<186> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[372] WL[373] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<187> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[374] WL[375] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<188> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[376] WL[377] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<189> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[378] WL[379] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<190> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[380] WL[381] S1AHSF400W40_MCB_2X4_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    MCB_508X4_SB_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_508X4_SB_CHAR BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] 
+ VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] 
+ WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] 
+ WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] 
+ WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] 
+ WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] 
+ WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] WL[64] WL[65] 
+ WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] 
+ WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] 
+ WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] 
+ WL[99] WL[100] WL[101] WL[102] WL[103] WL[104] WL[105] WL[106] WL[107] 
+ WL[108] WL[109] WL[110] WL[111] WL[112] WL[113] WL[114] WL[115] WL[116] 
+ WL[117] WL[118] WL[119] WL[120] WL[121] WL[122] WL[123] WL[124] WL[125] 
+ WL[126] WL[127] WL[128] WL[129] WL[130] WL[131] WL[132] WL[133] WL[134] 
+ WL[135] WL[136] WL[137] WL[138] WL[139] WL[140] WL[141] WL[142] WL[143] 
+ WL[144] WL[145] WL[146] WL[147] WL[148] WL[149] WL[150] WL[151] WL[152] 
+ WL[153] WL[154] WL[155] WL[156] WL[157] WL[158] WL[159] WL[160] WL[161] 
+ WL[162] WL[163] WL[164] WL[165] WL[166] WL[167] WL[168] WL[169] WL[170] 
+ WL[171] WL[172] WL[173] WL[174] WL[175] WL[176] WL[177] WL[178] WL[179] 
+ WL[180] WL[181] WL[182] WL[183] WL[184] WL[185] WL[186] WL[187] WL[188] 
+ WL[189] WL[190] WL[191] WL[192] WL[193] WL[194] WL[195] WL[196] WL[197] 
+ WL[198] WL[199] WL[200] WL[201] WL[202] WL[203] WL[204] WL[205] WL[206] 
+ WL[207] WL[208] WL[209] WL[210] WL[211] WL[212] WL[213] WL[214] WL[215] 
+ WL[216] WL[217] WL[218] WL[219] WL[220] WL[221] WL[222] WL[223] WL[224] 
+ WL[225] WL[226] WL[227] WL[228] WL[229] WL[230] WL[231] WL[232] WL[233] 
+ WL[234] WL[235] WL[236] WL[237] WL[238] WL[239] WL[240] WL[241] WL[242] 
+ WL[243] WL[244] WL[245] WL[246] WL[247] WL[248] WL[249] WL[250] WL[251] 
+ WL[252] WL[253] WL[254] WL[255] WL[256] WL[257] WL[258] WL[259] WL[260] 
+ WL[261] WL[262] WL[263] WL[264] WL[265] WL[266] WL[267] WL[268] WL[269] 
+ WL[270] WL[271] WL[272] WL[273] WL[274] WL[275] WL[276] WL[277] WL[278] 
+ WL[279] WL[280] WL[281] WL[282] WL[283] WL[284] WL[285] WL[286] WL[287] 
+ WL[288] WL[289] WL[290] WL[291] WL[292] WL[293] WL[294] WL[295] WL[296] 
+ WL[297] WL[298] WL[299] WL[300] WL[301] WL[302] WL[303] WL[304] WL[305] 
+ WL[306] WL[307] WL[308] WL[309] WL[310] WL[311] WL[312] WL[313] WL[314] 
+ WL[315] WL[316] WL[317] WL[318] WL[319] WL[320] WL[321] WL[322] WL[323] 
+ WL[324] WL[325] WL[326] WL[327] WL[328] WL[329] WL[330] WL[331] WL[332] 
+ WL[333] WL[334] WL[335] WL[336] WL[337] WL[338] WL[339] WL[340] WL[341] 
+ WL[342] WL[343] WL[344] WL[345] WL[346] WL[347] WL[348] WL[349] WL[350] 
+ WL[351] WL[352] WL[353] WL[354] WL[355] WL[356] WL[357] WL[358] WL[359] 
+ WL[360] WL[361] WL[362] WL[363] WL[364] WL[365] WL[366] WL[367] WL[368] 
+ WL[369] WL[370] WL[371] WL[372] WL[373] WL[374] WL[375] WL[376] WL[377] 
+ WL[378] WL[379] WL[380] WL[381] WL[382] WL[383] WL[384] WL[385] WL[386] 
+ WL[387] WL[388] WL[389] WL[390] WL[391] WL[392] WL[393] WL[394] WL[395] 
+ WL[396] WL[397] WL[398] WL[399] WL[400] WL[401] WL[402] WL[403] WL[404] 
+ WL[405] WL[406] WL[407] WL[408] WL[409] WL[410] WL[411] WL[412] WL[413] 
+ WL[414] WL[415] WL[416] WL[417] WL[418] WL[419] WL[420] WL[421] WL[422] 
+ WL[423] WL[424] WL[425] WL[426] WL[427] WL[428] WL[429] WL[430] WL[431] 
+ WL[432] WL[433] WL[434] WL[435] WL[436] WL[437] WL[438] WL[439] WL[440] 
+ WL[441] WL[442] WL[443] WL[444] WL[445] WL[446] WL[447] WL[448] WL[449] 
+ WL[450] WL[451] WL[452] WL[453] WL[454] WL[455] WL[456] WL[457] WL[458] 
+ WL[459] WL[460] WL[461] WL[462] WL[463] WL[464] WL[465] WL[466] WL[467] 
+ WL[468] WL[469] WL[470] WL[471] WL[472] WL[473] WL[474] WL[475] WL[476] 
+ WL[477] WL[478] WL[479] WL[480] WL[481] WL[482] WL[483] WL[484] WL[485] 
+ WL[486] WL[487] WL[488] WL[489] WL[490] WL[491] WL[492] WL[493] WL[494] 
+ WL[495] WL[496] WL[497] WL[498] WL[499] WL[500] WL[501] WL[502] WL[503] 
+ WL[504] WL[505] WL[506] WL[507]
*.PININFO WL[0]:I WL[1]:I WL[2]:I WL[3]:I WL[4]:I WL[5]:I WL[6]:I WL[7]:I 
*.PININFO WL[8]:I WL[9]:I WL[10]:I WL[11]:I WL[12]:I WL[13]:I WL[14]:I 
*.PININFO WL[15]:I WL[16]:I WL[17]:I WL[18]:I WL[19]:I WL[20]:I WL[21]:I 
*.PININFO WL[22]:I WL[23]:I WL[24]:I WL[25]:I WL[26]:I WL[27]:I WL[28]:I 
*.PININFO WL[29]:I WL[30]:I WL[31]:I WL[32]:I WL[33]:I WL[34]:I WL[35]:I 
*.PININFO WL[36]:I WL[37]:I WL[38]:I WL[39]:I WL[40]:I WL[41]:I WL[42]:I 
*.PININFO WL[43]:I WL[44]:I WL[45]:I WL[46]:I WL[47]:I WL[48]:I WL[49]:I 
*.PININFO WL[50]:I WL[51]:I WL[52]:I WL[53]:I WL[54]:I WL[55]:I WL[56]:I 
*.PININFO WL[57]:I WL[58]:I WL[59]:I WL[60]:I WL[61]:I WL[62]:I WL[63]:I 
*.PININFO WL[64]:I WL[65]:I WL[66]:I WL[67]:I WL[68]:I WL[69]:I WL[70]:I 
*.PININFO WL[71]:I WL[72]:I WL[73]:I WL[74]:I WL[75]:I WL[76]:I WL[77]:I 
*.PININFO WL[78]:I WL[79]:I WL[80]:I WL[81]:I WL[82]:I WL[83]:I WL[84]:I 
*.PININFO WL[85]:I WL[86]:I WL[87]:I WL[88]:I WL[89]:I WL[90]:I WL[91]:I 
*.PININFO WL[92]:I WL[93]:I WL[94]:I WL[95]:I WL[96]:I WL[97]:I WL[98]:I 
*.PININFO WL[99]:I WL[100]:I WL[101]:I WL[102]:I WL[103]:I WL[104]:I WL[105]:I 
*.PININFO WL[106]:I WL[107]:I WL[108]:I WL[109]:I WL[110]:I WL[111]:I 
*.PININFO WL[112]:I WL[113]:I WL[114]:I WL[115]:I WL[116]:I WL[117]:I 
*.PININFO WL[118]:I WL[119]:I WL[120]:I WL[121]:I WL[122]:I WL[123]:I 
*.PININFO WL[124]:I WL[125]:I WL[126]:I WL[127]:I WL[128]:I WL[129]:I 
*.PININFO WL[130]:I WL[131]:I WL[132]:I WL[133]:I WL[134]:I WL[135]:I 
*.PININFO WL[136]:I WL[137]:I WL[138]:I WL[139]:I WL[140]:I WL[141]:I 
*.PININFO WL[142]:I WL[143]:I WL[144]:I WL[145]:I WL[146]:I WL[147]:I 
*.PININFO WL[148]:I WL[149]:I WL[150]:I WL[151]:I WL[152]:I WL[153]:I 
*.PININFO WL[154]:I WL[155]:I WL[156]:I WL[157]:I WL[158]:I WL[159]:I 
*.PININFO WL[160]:I WL[161]:I WL[162]:I WL[163]:I WL[164]:I WL[165]:I 
*.PININFO WL[166]:I WL[167]:I WL[168]:I WL[169]:I WL[170]:I WL[171]:I 
*.PININFO WL[172]:I WL[173]:I WL[174]:I WL[175]:I WL[176]:I WL[177]:I 
*.PININFO WL[178]:I WL[179]:I WL[180]:I WL[181]:I WL[182]:I WL[183]:I 
*.PININFO WL[184]:I WL[185]:I WL[186]:I WL[187]:I WL[188]:I WL[189]:I 
*.PININFO WL[190]:I WL[191]:I WL[192]:I WL[193]:I WL[194]:I WL[195]:I 
*.PININFO WL[196]:I WL[197]:I WL[198]:I WL[199]:I WL[200]:I WL[201]:I 
*.PININFO WL[202]:I WL[203]:I WL[204]:I WL[205]:I WL[206]:I WL[207]:I 
*.PININFO WL[208]:I WL[209]:I WL[210]:I WL[211]:I WL[212]:I WL[213]:I 
*.PININFO WL[214]:I WL[215]:I WL[216]:I WL[217]:I WL[218]:I WL[219]:I 
*.PININFO WL[220]:I WL[221]:I WL[222]:I WL[223]:I WL[224]:I WL[225]:I 
*.PININFO WL[226]:I WL[227]:I WL[228]:I WL[229]:I WL[230]:I WL[231]:I 
*.PININFO WL[232]:I WL[233]:I WL[234]:I WL[235]:I WL[236]:I WL[237]:I 
*.PININFO WL[238]:I WL[239]:I WL[240]:I WL[241]:I WL[242]:I WL[243]:I 
*.PININFO WL[244]:I WL[245]:I WL[246]:I WL[247]:I WL[248]:I WL[249]:I 
*.PININFO WL[250]:I WL[251]:I WL[252]:I WL[253]:I WL[254]:I WL[255]:I 
*.PININFO WL[256]:I WL[257]:I WL[258]:I WL[259]:I WL[260]:I WL[261]:I 
*.PININFO WL[262]:I WL[263]:I WL[264]:I WL[265]:I WL[266]:I WL[267]:I 
*.PININFO WL[268]:I WL[269]:I WL[270]:I WL[271]:I WL[272]:I WL[273]:I 
*.PININFO WL[274]:I WL[275]:I WL[276]:I WL[277]:I WL[278]:I WL[279]:I 
*.PININFO WL[280]:I WL[281]:I WL[282]:I WL[283]:I WL[284]:I WL[285]:I 
*.PININFO WL[286]:I WL[287]:I WL[288]:I WL[289]:I WL[290]:I WL[291]:I 
*.PININFO WL[292]:I WL[293]:I WL[294]:I WL[295]:I WL[296]:I WL[297]:I 
*.PININFO WL[298]:I WL[299]:I WL[300]:I WL[301]:I WL[302]:I WL[303]:I 
*.PININFO WL[304]:I WL[305]:I WL[306]:I WL[307]:I WL[308]:I WL[309]:I 
*.PININFO WL[310]:I WL[311]:I WL[312]:I WL[313]:I WL[314]:I WL[315]:I 
*.PININFO WL[316]:I WL[317]:I WL[318]:I WL[319]:I WL[320]:I WL[321]:I 
*.PININFO WL[322]:I WL[323]:I WL[324]:I WL[325]:I WL[326]:I WL[327]:I 
*.PININFO WL[328]:I WL[329]:I WL[330]:I WL[331]:I WL[332]:I WL[333]:I 
*.PININFO WL[334]:I WL[335]:I WL[336]:I WL[337]:I WL[338]:I WL[339]:I 
*.PININFO WL[340]:I WL[341]:I WL[342]:I WL[343]:I WL[344]:I WL[345]:I 
*.PININFO WL[346]:I WL[347]:I WL[348]:I WL[349]:I WL[350]:I WL[351]:I 
*.PININFO WL[352]:I WL[353]:I WL[354]:I WL[355]:I WL[356]:I WL[357]:I 
*.PININFO WL[358]:I WL[359]:I WL[360]:I WL[361]:I WL[362]:I WL[363]:I 
*.PININFO WL[364]:I WL[365]:I WL[366]:I WL[367]:I WL[368]:I WL[369]:I 
*.PININFO WL[370]:I WL[371]:I WL[372]:I WL[373]:I WL[374]:I WL[375]:I 
*.PININFO WL[376]:I WL[377]:I WL[378]:I WL[379]:I WL[380]:I WL[381]:I 
*.PININFO WL[382]:I WL[383]:I WL[384]:I WL[385]:I WL[386]:I WL[387]:I 
*.PININFO WL[388]:I WL[389]:I WL[390]:I WL[391]:I WL[392]:I WL[393]:I 
*.PININFO WL[394]:I WL[395]:I WL[396]:I WL[397]:I WL[398]:I WL[399]:I 
*.PININFO WL[400]:I WL[401]:I WL[402]:I WL[403]:I WL[404]:I WL[405]:I 
*.PININFO WL[406]:I WL[407]:I WL[408]:I WL[409]:I WL[410]:I WL[411]:I 
*.PININFO WL[412]:I WL[413]:I WL[414]:I WL[415]:I WL[416]:I WL[417]:I 
*.PININFO WL[418]:I WL[419]:I WL[420]:I WL[421]:I WL[422]:I WL[423]:I 
*.PININFO WL[424]:I WL[425]:I WL[426]:I WL[427]:I WL[428]:I WL[429]:I 
*.PININFO WL[430]:I WL[431]:I WL[432]:I WL[433]:I WL[434]:I WL[435]:I 
*.PININFO WL[436]:I WL[437]:I WL[438]:I WL[439]:I WL[440]:I WL[441]:I 
*.PININFO WL[442]:I WL[443]:I WL[444]:I WL[445]:I WL[446]:I WL[447]:I 
*.PININFO WL[448]:I WL[449]:I WL[450]:I WL[451]:I WL[452]:I WL[453]:I 
*.PININFO WL[454]:I WL[455]:I WL[456]:I WL[457]:I WL[458]:I WL[459]:I 
*.PININFO WL[460]:I WL[461]:I WL[462]:I WL[463]:I WL[464]:I WL[465]:I 
*.PININFO WL[466]:I WL[467]:I WL[468]:I WL[469]:I WL[470]:I WL[471]:I 
*.PININFO WL[472]:I WL[473]:I WL[474]:I WL[475]:I WL[476]:I WL[477]:I 
*.PININFO WL[478]:I WL[479]:I WL[480]:I WL[481]:I WL[482]:I WL[483]:I 
*.PININFO WL[484]:I WL[485]:I WL[486]:I WL[487]:I WL[488]:I WL[489]:I 
*.PININFO WL[490]:I WL[491]:I WL[492]:I WL[493]:I WL[494]:I WL[495]:I 
*.PININFO WL[496]:I WL[497]:I WL[498]:I WL[499]:I WL[500]:I WL[501]:I 
*.PININFO WL[502]:I WL[503]:I WL[504]:I WL[505]:I WL[506]:I WL[507]:I BL[0]:B 
*.PININFO BL[1]:B BL[2]:B BL[3]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B VDDI:B 
*.PININFO VSSI:B
XMCB_2X4<0> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[0] WL[1] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<1> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[2] WL[3] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<2> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[4] WL[5] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<3> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[6] WL[7] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<4> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[8] WL[9] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<5> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[10] WL[11] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<6> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[12] WL[13] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<7> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[14] WL[15] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<8> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[16] WL[17] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<9> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[18] WL[19] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<10> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[20] WL[21] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<11> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[22] WL[23] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<12> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[24] WL[25] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<13> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[26] WL[27] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<14> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[28] WL[29] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<15> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[30] WL[31] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<16> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[32] WL[33] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<17> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[34] WL[35] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<18> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[36] WL[37] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<19> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[38] WL[39] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<20> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[40] WL[41] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<21> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[42] WL[43] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<22> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[44] WL[45] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<23> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[46] WL[47] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<24> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[48] WL[49] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<25> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[50] WL[51] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<26> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[52] WL[53] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<27> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[54] WL[55] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<28> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[56] WL[57] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<29> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[58] WL[59] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<30> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[60] WL[61] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<31> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[62] WL[63] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<32> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[64] WL[65] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<33> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[66] WL[67] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<34> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[68] WL[69] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<35> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[70] WL[71] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<36> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[72] WL[73] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<37> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[74] WL[75] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<38> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[76] WL[77] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<39> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[78] WL[79] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<40> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[80] WL[81] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<41> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[82] WL[83] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<42> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[84] WL[85] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<43> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[86] WL[87] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<44> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[88] WL[89] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<45> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[90] WL[91] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<46> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[92] WL[93] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<47> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[94] WL[95] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<48> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[96] WL[97] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<49> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[98] WL[99] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<50> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[100] WL[101] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<51> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[102] WL[103] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<52> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[104] WL[105] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<53> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[106] WL[107] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<54> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[108] WL[109] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<55> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[110] WL[111] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<56> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[112] WL[113] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<57> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[114] WL[115] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<58> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[116] WL[117] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<59> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[118] WL[119] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<60> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[120] WL[121] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<61> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[122] WL[123] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<62> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[124] WL[125] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<63> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[126] WL[127] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<64> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[128] WL[129] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<65> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[130] WL[131] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<66> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[132] WL[133] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<67> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[134] WL[135] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<68> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[136] WL[137] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<69> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[138] WL[139] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<70> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[140] WL[141] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<71> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[142] WL[143] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<72> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[144] WL[145] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<73> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[146] WL[147] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<74> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[148] WL[149] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<75> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[150] WL[151] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<76> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[152] WL[153] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<77> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[154] WL[155] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<78> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[156] WL[157] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<79> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[158] WL[159] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<80> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[160] WL[161] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<81> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[162] WL[163] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<82> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[164] WL[165] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<83> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[166] WL[167] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<84> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[168] WL[169] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<85> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[170] WL[171] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<86> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[172] WL[173] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<87> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[174] WL[175] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<88> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[176] WL[177] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<89> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[178] WL[179] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<90> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[180] WL[181] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<91> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[182] WL[183] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<92> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[184] WL[185] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<93> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[186] WL[187] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<94> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[188] WL[189] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<95> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[190] WL[191] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<96> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[192] WL[193] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<97> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[194] WL[195] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<98> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[196] WL[197] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<99> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[198] WL[199] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<100> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[200] WL[201] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<101> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[202] WL[203] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<102> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[204] WL[205] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<103> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[206] WL[207] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<104> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[208] WL[209] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<105> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[210] WL[211] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<106> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[212] WL[213] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<107> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[214] WL[215] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<108> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[216] WL[217] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<109> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[218] WL[219] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<110> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[220] WL[221] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<111> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[222] WL[223] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<112> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[224] WL[225] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<113> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[226] WL[227] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<114> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[228] WL[229] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<115> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[230] WL[231] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<116> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[232] WL[233] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<117> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[234] WL[235] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<118> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[236] WL[237] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<119> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[238] WL[239] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<120> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[240] WL[241] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<121> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[242] WL[243] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<122> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[244] WL[245] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<123> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[246] WL[247] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<124> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[248] WL[249] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<125> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[250] WL[251] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<126> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[252] WL[253] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<127> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[254] WL[255] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<128> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[256] WL[257] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<129> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[258] WL[259] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<130> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[260] WL[261] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<131> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[262] WL[263] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<132> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[264] WL[265] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<133> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[266] WL[267] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<134> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[268] WL[269] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<135> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[270] WL[271] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<136> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[272] WL[273] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<137> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[274] WL[275] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<138> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[276] WL[277] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<139> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[278] WL[279] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<140> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[280] WL[281] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<141> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[282] WL[283] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<142> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[284] WL[285] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<143> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[286] WL[287] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<144> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[288] WL[289] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<145> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[290] WL[291] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<146> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[292] WL[293] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<147> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[294] WL[295] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<148> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[296] WL[297] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<149> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[298] WL[299] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<150> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[300] WL[301] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<151> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[302] WL[303] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<152> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[304] WL[305] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<153> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[306] WL[307] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<154> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[308] WL[309] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<155> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[310] WL[311] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<156> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[312] WL[313] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<157> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[314] WL[315] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<158> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[316] WL[317] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<159> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[318] WL[319] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<160> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[320] WL[321] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<161> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[322] WL[323] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<162> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[324] WL[325] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<163> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[326] WL[327] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<164> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[328] WL[329] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<165> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[330] WL[331] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<166> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[332] WL[333] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<167> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[334] WL[335] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<168> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[336] WL[337] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<169> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[338] WL[339] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<170> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[340] WL[341] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<171> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[342] WL[343] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<172> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[344] WL[345] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<173> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[346] WL[347] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<174> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[348] WL[349] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<175> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[350] WL[351] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<176> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[352] WL[353] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<177> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[354] WL[355] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<178> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[356] WL[357] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<179> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[358] WL[359] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<180> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[360] WL[361] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<181> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[362] WL[363] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<182> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[364] WL[365] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<183> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[366] WL[367] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<184> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[368] WL[369] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<185> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[370] WL[371] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<186> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[372] WL[373] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<187> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[374] WL[375] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<188> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[376] WL[377] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<189> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[378] WL[379] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<190> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[380] WL[381] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<191> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[382] WL[383] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<192> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[384] WL[385] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<193> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[386] WL[387] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<194> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[388] WL[389] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<195> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[390] WL[391] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<196> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[392] WL[393] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<197> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[394] WL[395] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<198> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[396] WL[397] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<199> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[398] WL[399] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<200> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[400] WL[401] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<201> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[402] WL[403] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<202> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[404] WL[405] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<203> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[406] WL[407] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<204> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[408] WL[409] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<205> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[410] WL[411] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<206> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[412] WL[413] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<207> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[414] WL[415] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<208> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[416] WL[417] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<209> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[418] WL[419] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<210> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[420] WL[421] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<211> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[422] WL[423] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<212> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[424] WL[425] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<213> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[426] WL[427] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<214> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[428] WL[429] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<215> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[430] WL[431] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<216> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[432] WL[433] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<217> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[434] WL[435] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<218> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[436] WL[437] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<219> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[438] WL[439] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<220> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[440] WL[441] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<221> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[442] WL[443] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<222> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[444] WL[445] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<223> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[446] WL[447] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<224> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[448] WL[449] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<225> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[450] WL[451] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<226> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[452] WL[453] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<227> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[454] WL[455] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<228> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[456] WL[457] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<229> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[458] WL[459] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<230> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[460] WL[461] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<231> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[462] WL[463] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<232> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[464] WL[465] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<233> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[466] WL[467] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<234> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[468] WL[469] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<235> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[470] WL[471] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<236> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[472] WL[473] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<237> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[474] WL[475] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<238> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[476] WL[477] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<239> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[478] WL[479] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<240> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[480] WL[481] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<241> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[482] WL[483] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<242> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[484] WL[485] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<243> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[486] WL[487] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<244> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[488] WL[489] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<245> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[490] WL[491] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<246> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[492] WL[493] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<247> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[494] WL[495] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<248> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[496] WL[497] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<249> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[498] WL[499] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<250> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[500] WL[501] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<251> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[502] WL[503] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<252> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[504] WL[505] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<253> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[506] WL[507] S1AHSF400W40_MCB_2X4_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    MCB_254X4_SB_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_254X4_SB_CHAR BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] 
+ VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] 
+ WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] 
+ WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] 
+ WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] 
+ WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] 
+ WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] WL[64] WL[65] 
+ WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] 
+ WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] 
+ WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] 
+ WL[99] WL[100] WL[101] WL[102] WL[103] WL[104] WL[105] WL[106] WL[107] 
+ WL[108] WL[109] WL[110] WL[111] WL[112] WL[113] WL[114] WL[115] WL[116] 
+ WL[117] WL[118] WL[119] WL[120] WL[121] WL[122] WL[123] WL[124] WL[125] 
+ WL[126] WL[127] WL[128] WL[129] WL[130] WL[131] WL[132] WL[133] WL[134] 
+ WL[135] WL[136] WL[137] WL[138] WL[139] WL[140] WL[141] WL[142] WL[143] 
+ WL[144] WL[145] WL[146] WL[147] WL[148] WL[149] WL[150] WL[151] WL[152] 
+ WL[153] WL[154] WL[155] WL[156] WL[157] WL[158] WL[159] WL[160] WL[161] 
+ WL[162] WL[163] WL[164] WL[165] WL[166] WL[167] WL[168] WL[169] WL[170] 
+ WL[171] WL[172] WL[173] WL[174] WL[175] WL[176] WL[177] WL[178] WL[179] 
+ WL[180] WL[181] WL[182] WL[183] WL[184] WL[185] WL[186] WL[187] WL[188] 
+ WL[189] WL[190] WL[191] WL[192] WL[193] WL[194] WL[195] WL[196] WL[197] 
+ WL[198] WL[199] WL[200] WL[201] WL[202] WL[203] WL[204] WL[205] WL[206] 
+ WL[207] WL[208] WL[209] WL[210] WL[211] WL[212] WL[213] WL[214] WL[215] 
+ WL[216] WL[217] WL[218] WL[219] WL[220] WL[221] WL[222] WL[223] WL[224] 
+ WL[225] WL[226] WL[227] WL[228] WL[229] WL[230] WL[231] WL[232] WL[233] 
+ WL[234] WL[235] WL[236] WL[237] WL[238] WL[239] WL[240] WL[241] WL[242] 
+ WL[243] WL[244] WL[245] WL[246] WL[247] WL[248] WL[249] WL[250] WL[251] 
+ WL[252] WL[253]
*.PININFO WL[0]:I WL[1]:I WL[2]:I WL[3]:I WL[4]:I WL[5]:I WL[6]:I WL[7]:I 
*.PININFO WL[8]:I WL[9]:I WL[10]:I WL[11]:I WL[12]:I WL[13]:I WL[14]:I 
*.PININFO WL[15]:I WL[16]:I WL[17]:I WL[18]:I WL[19]:I WL[20]:I WL[21]:I 
*.PININFO WL[22]:I WL[23]:I WL[24]:I WL[25]:I WL[26]:I WL[27]:I WL[28]:I 
*.PININFO WL[29]:I WL[30]:I WL[31]:I WL[32]:I WL[33]:I WL[34]:I WL[35]:I 
*.PININFO WL[36]:I WL[37]:I WL[38]:I WL[39]:I WL[40]:I WL[41]:I WL[42]:I 
*.PININFO WL[43]:I WL[44]:I WL[45]:I WL[46]:I WL[47]:I WL[48]:I WL[49]:I 
*.PININFO WL[50]:I WL[51]:I WL[52]:I WL[53]:I WL[54]:I WL[55]:I WL[56]:I 
*.PININFO WL[57]:I WL[58]:I WL[59]:I WL[60]:I WL[61]:I WL[62]:I WL[63]:I 
*.PININFO WL[64]:I WL[65]:I WL[66]:I WL[67]:I WL[68]:I WL[69]:I WL[70]:I 
*.PININFO WL[71]:I WL[72]:I WL[73]:I WL[74]:I WL[75]:I WL[76]:I WL[77]:I 
*.PININFO WL[78]:I WL[79]:I WL[80]:I WL[81]:I WL[82]:I WL[83]:I WL[84]:I 
*.PININFO WL[85]:I WL[86]:I WL[87]:I WL[88]:I WL[89]:I WL[90]:I WL[91]:I 
*.PININFO WL[92]:I WL[93]:I WL[94]:I WL[95]:I WL[96]:I WL[97]:I WL[98]:I 
*.PININFO WL[99]:I WL[100]:I WL[101]:I WL[102]:I WL[103]:I WL[104]:I WL[105]:I 
*.PININFO WL[106]:I WL[107]:I WL[108]:I WL[109]:I WL[110]:I WL[111]:I 
*.PININFO WL[112]:I WL[113]:I WL[114]:I WL[115]:I WL[116]:I WL[117]:I 
*.PININFO WL[118]:I WL[119]:I WL[120]:I WL[121]:I WL[122]:I WL[123]:I 
*.PININFO WL[124]:I WL[125]:I WL[126]:I WL[127]:I WL[128]:I WL[129]:I 
*.PININFO WL[130]:I WL[131]:I WL[132]:I WL[133]:I WL[134]:I WL[135]:I 
*.PININFO WL[136]:I WL[137]:I WL[138]:I WL[139]:I WL[140]:I WL[141]:I 
*.PININFO WL[142]:I WL[143]:I WL[144]:I WL[145]:I WL[146]:I WL[147]:I 
*.PININFO WL[148]:I WL[149]:I WL[150]:I WL[151]:I WL[152]:I WL[153]:I 
*.PININFO WL[154]:I WL[155]:I WL[156]:I WL[157]:I WL[158]:I WL[159]:I 
*.PININFO WL[160]:I WL[161]:I WL[162]:I WL[163]:I WL[164]:I WL[165]:I 
*.PININFO WL[166]:I WL[167]:I WL[168]:I WL[169]:I WL[170]:I WL[171]:I 
*.PININFO WL[172]:I WL[173]:I WL[174]:I WL[175]:I WL[176]:I WL[177]:I 
*.PININFO WL[178]:I WL[179]:I WL[180]:I WL[181]:I WL[182]:I WL[183]:I 
*.PININFO WL[184]:I WL[185]:I WL[186]:I WL[187]:I WL[188]:I WL[189]:I 
*.PININFO WL[190]:I WL[191]:I WL[192]:I WL[193]:I WL[194]:I WL[195]:I 
*.PININFO WL[196]:I WL[197]:I WL[198]:I WL[199]:I WL[200]:I WL[201]:I 
*.PININFO WL[202]:I WL[203]:I WL[204]:I WL[205]:I WL[206]:I WL[207]:I 
*.PININFO WL[208]:I WL[209]:I WL[210]:I WL[211]:I WL[212]:I WL[213]:I 
*.PININFO WL[214]:I WL[215]:I WL[216]:I WL[217]:I WL[218]:I WL[219]:I 
*.PININFO WL[220]:I WL[221]:I WL[222]:I WL[223]:I WL[224]:I WL[225]:I 
*.PININFO WL[226]:I WL[227]:I WL[228]:I WL[229]:I WL[230]:I WL[231]:I 
*.PININFO WL[232]:I WL[233]:I WL[234]:I WL[235]:I WL[236]:I WL[237]:I 
*.PININFO WL[238]:I WL[239]:I WL[240]:I WL[241]:I WL[242]:I WL[243]:I 
*.PININFO WL[244]:I WL[245]:I WL[246]:I WL[247]:I WL[248]:I WL[249]:I 
*.PININFO WL[250]:I WL[251]:I WL[252]:I WL[253]:I BL[0]:B BL[1]:B BL[2]:B 
*.PININFO BL[3]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B VDDI:B VSSI:B
XMCB_2X4<0> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[0] WL[1] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<1> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[2] WL[3] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<2> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[4] WL[5] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<3> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[6] WL[7] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<4> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[8] WL[9] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<5> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[10] WL[11] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<6> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[12] WL[13] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<7> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[14] WL[15] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<8> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[16] WL[17] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<9> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[18] WL[19] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<10> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[20] WL[21] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<11> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[22] WL[23] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<12> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[24] WL[25] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<13> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[26] WL[27] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<14> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[28] WL[29] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<15> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[30] WL[31] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<16> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[32] WL[33] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<17> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[34] WL[35] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<18> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[36] WL[37] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<19> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[38] WL[39] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<20> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[40] WL[41] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<21> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[42] WL[43] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<22> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[44] WL[45] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<23> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[46] WL[47] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<24> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[48] WL[49] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<25> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[50] WL[51] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<26> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[52] WL[53] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<27> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[54] WL[55] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<28> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[56] WL[57] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<29> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[58] WL[59] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<30> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[60] WL[61] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<31> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[62] WL[63] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<32> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[64] WL[65] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<33> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[66] WL[67] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<34> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[68] WL[69] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<35> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[70] WL[71] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<36> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[72] WL[73] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<37> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[74] WL[75] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<38> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[76] WL[77] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<39> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[78] WL[79] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<40> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[80] WL[81] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<41> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[82] WL[83] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<42> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[84] WL[85] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<43> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[86] WL[87] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<44> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[88] WL[89] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<45> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[90] WL[91] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<46> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[92] WL[93] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<47> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[94] WL[95] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<48> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[96] WL[97] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<49> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[98] WL[99] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<50> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[100] WL[101] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<51> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[102] WL[103] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<52> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[104] WL[105] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<53> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[106] WL[107] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<54> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[108] WL[109] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<55> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[110] WL[111] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<56> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[112] WL[113] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<57> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[114] WL[115] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<58> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[116] WL[117] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<59> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[118] WL[119] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<60> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[120] WL[121] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<61> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[122] WL[123] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<62> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[124] WL[125] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<63> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[126] WL[127] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<64> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[128] WL[129] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<65> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[130] WL[131] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<66> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[132] WL[133] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<67> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[134] WL[135] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<68> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[136] WL[137] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<69> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[138] WL[139] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<70> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[140] WL[141] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<71> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[142] WL[143] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<72> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[144] WL[145] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<73> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[146] WL[147] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<74> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[148] WL[149] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<75> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[150] WL[151] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<76> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[152] WL[153] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<77> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[154] WL[155] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<78> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[156] WL[157] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<79> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[158] WL[159] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<80> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[160] WL[161] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<81> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[162] WL[163] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<82> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[164] WL[165] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<83> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[166] WL[167] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<84> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[168] WL[169] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<85> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[170] WL[171] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<86> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[172] WL[173] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<87> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[174] WL[175] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<88> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[176] WL[177] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<89> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[178] WL[179] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<90> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[180] WL[181] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<91> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[182] WL[183] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<92> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[184] WL[185] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<93> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[186] WL[187] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<94> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[188] WL[189] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<95> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[190] WL[191] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<96> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[192] WL[193] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<97> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[194] WL[195] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<98> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[196] WL[197] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<99> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[198] WL[199] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<100> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[200] WL[201] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<101> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[202] WL[203] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<102> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[204] WL[205] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<103> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[206] WL[207] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<104> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[208] WL[209] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<105> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[210] WL[211] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<106> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[212] WL[213] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<107> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[214] WL[215] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<108> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[216] WL[217] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<109> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[218] WL[219] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<110> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[220] WL[221] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<111> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[222] WL[223] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<112> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[224] WL[225] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<113> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[226] WL[227] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<114> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[228] WL[229] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<115> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[230] WL[231] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<116> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[232] WL[233] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<117> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[234] WL[235] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<118> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[236] WL[237] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<119> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[238] WL[239] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<120> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[240] WL[241] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<121> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[242] WL[243] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<122> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[244] WL[245] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<123> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[246] WL[247] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<124> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[248] WL[249] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<125> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[250] WL[251] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<126> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[252] WL[253] S1AHSF400W40_MCB_2X4_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    MCB_126X4_SB_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_126X4_SB_CHAR BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] 
+ VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] 
+ WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] 
+ WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] 
+ WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] 
+ WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] 
+ WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] WL[64] WL[65] 
+ WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] 
+ WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] 
+ WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] 
+ WL[99] WL[100] WL[101] WL[102] WL[103] WL[104] WL[105] WL[106] WL[107] 
+ WL[108] WL[109] WL[110] WL[111] WL[112] WL[113] WL[114] WL[115] WL[116] 
+ WL[117] WL[118] WL[119] WL[120] WL[121] WL[122] WL[123] WL[124] WL[125]
*.PININFO WL[0]:I WL[1]:I WL[2]:I WL[3]:I WL[4]:I WL[5]:I WL[6]:I WL[7]:I 
*.PININFO WL[8]:I WL[9]:I WL[10]:I WL[11]:I WL[12]:I WL[13]:I WL[14]:I 
*.PININFO WL[15]:I WL[16]:I WL[17]:I WL[18]:I WL[19]:I WL[20]:I WL[21]:I 
*.PININFO WL[22]:I WL[23]:I WL[24]:I WL[25]:I WL[26]:I WL[27]:I WL[28]:I 
*.PININFO WL[29]:I WL[30]:I WL[31]:I WL[32]:I WL[33]:I WL[34]:I WL[35]:I 
*.PININFO WL[36]:I WL[37]:I WL[38]:I WL[39]:I WL[40]:I WL[41]:I WL[42]:I 
*.PININFO WL[43]:I WL[44]:I WL[45]:I WL[46]:I WL[47]:I WL[48]:I WL[49]:I 
*.PININFO WL[50]:I WL[51]:I WL[52]:I WL[53]:I WL[54]:I WL[55]:I WL[56]:I 
*.PININFO WL[57]:I WL[58]:I WL[59]:I WL[60]:I WL[61]:I WL[62]:I WL[63]:I 
*.PININFO WL[64]:I WL[65]:I WL[66]:I WL[67]:I WL[68]:I WL[69]:I WL[70]:I 
*.PININFO WL[71]:I WL[72]:I WL[73]:I WL[74]:I WL[75]:I WL[76]:I WL[77]:I 
*.PININFO WL[78]:I WL[79]:I WL[80]:I WL[81]:I WL[82]:I WL[83]:I WL[84]:I 
*.PININFO WL[85]:I WL[86]:I WL[87]:I WL[88]:I WL[89]:I WL[90]:I WL[91]:I 
*.PININFO WL[92]:I WL[93]:I WL[94]:I WL[95]:I WL[96]:I WL[97]:I WL[98]:I 
*.PININFO WL[99]:I WL[100]:I WL[101]:I WL[102]:I WL[103]:I WL[104]:I WL[105]:I 
*.PININFO WL[106]:I WL[107]:I WL[108]:I WL[109]:I WL[110]:I WL[111]:I 
*.PININFO WL[112]:I WL[113]:I WL[114]:I WL[115]:I WL[116]:I WL[117]:I 
*.PININFO WL[118]:I WL[119]:I WL[120]:I WL[121]:I WL[122]:I WL[123]:I 
*.PININFO WL[124]:I WL[125]:I BL[0]:B BL[1]:B BL[2]:B BL[3]:B BLB[0]:B 
*.PININFO BLB[1]:B BLB[2]:B BLB[3]:B VDDI:B VSSI:B
XMCB_2X4<0> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[0] WL[1] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<1> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[2] WL[3] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<2> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[4] WL[5] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<3> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[6] WL[7] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<4> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[8] WL[9] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<5> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[10] WL[11] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<6> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[12] WL[13] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<7> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[14] WL[15] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<8> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[16] WL[17] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<9> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[18] WL[19] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<10> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[20] WL[21] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<11> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[22] WL[23] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<12> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[24] WL[25] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<13> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[26] WL[27] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<14> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[28] WL[29] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<15> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[30] WL[31] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<16> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[32] WL[33] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<17> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[34] WL[35] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<18> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[36] WL[37] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<19> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[38] WL[39] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<20> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[40] WL[41] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<21> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[42] WL[43] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<22> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[44] WL[45] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<23> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[46] WL[47] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<24> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[48] WL[49] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<25> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[50] WL[51] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<26> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[52] WL[53] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<27> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[54] WL[55] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<28> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[56] WL[57] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<29> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[58] WL[59] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<30> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[60] WL[61] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<31> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[62] WL[63] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<32> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[64] WL[65] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<33> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[66] WL[67] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<34> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[68] WL[69] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<35> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[70] WL[71] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<36> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[72] WL[73] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<37> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[74] WL[75] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<38> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[76] WL[77] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<39> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[78] WL[79] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<40> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[80] WL[81] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<41> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[82] WL[83] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<42> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[84] WL[85] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<43> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[86] WL[87] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<44> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[88] WL[89] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<45> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[90] WL[91] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<46> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[92] WL[93] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<47> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[94] WL[95] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<48> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[96] WL[97] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<49> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[98] WL[99] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<50> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[100] WL[101] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<51> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[102] WL[103] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<52> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[104] WL[105] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<53> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[106] WL[107] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<54> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[108] WL[109] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<55> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[110] WL[111] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<56> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[112] WL[113] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<57> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[114] WL[115] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<58> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[116] WL[117] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<59> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[118] WL[119] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<60> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[120] WL[121] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<61> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[122] WL[123] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<62> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[124] WL[125] S1AHSF400W40_MCB_2X4_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    MCB_252X4_SB_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_252X4_SB_CHAR BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] 
+ VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] 
+ WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] 
+ WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] 
+ WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] 
+ WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] 
+ WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] WL[64] WL[65] 
+ WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] 
+ WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] 
+ WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] 
+ WL[99] WL[100] WL[101] WL[102] WL[103] WL[104] WL[105] WL[106] WL[107] 
+ WL[108] WL[109] WL[110] WL[111] WL[112] WL[113] WL[114] WL[115] WL[116] 
+ WL[117] WL[118] WL[119] WL[120] WL[121] WL[122] WL[123] WL[124] WL[125] 
+ WL[126] WL[127] WL[128] WL[129] WL[130] WL[131] WL[132] WL[133] WL[134] 
+ WL[135] WL[136] WL[137] WL[138] WL[139] WL[140] WL[141] WL[142] WL[143] 
+ WL[144] WL[145] WL[146] WL[147] WL[148] WL[149] WL[150] WL[151] WL[152] 
+ WL[153] WL[154] WL[155] WL[156] WL[157] WL[158] WL[159] WL[160] WL[161] 
+ WL[162] WL[163] WL[164] WL[165] WL[166] WL[167] WL[168] WL[169] WL[170] 
+ WL[171] WL[172] WL[173] WL[174] WL[175] WL[176] WL[177] WL[178] WL[179] 
+ WL[180] WL[181] WL[182] WL[183] WL[184] WL[185] WL[186] WL[187] WL[188] 
+ WL[189] WL[190] WL[191] WL[192] WL[193] WL[194] WL[195] WL[196] WL[197] 
+ WL[198] WL[199] WL[200] WL[201] WL[202] WL[203] WL[204] WL[205] WL[206] 
+ WL[207] WL[208] WL[209] WL[210] WL[211] WL[212] WL[213] WL[214] WL[215] 
+ WL[216] WL[217] WL[218] WL[219] WL[220] WL[221] WL[222] WL[223] WL[224] 
+ WL[225] WL[226] WL[227] WL[228] WL[229] WL[230] WL[231] WL[232] WL[233] 
+ WL[234] WL[235] WL[236] WL[237] WL[238] WL[239] WL[240] WL[241] WL[242] 
+ WL[243] WL[244] WL[245] WL[246] WL[247] WL[248] WL[249] WL[250] WL[251]
*.PININFO WL[0]:I WL[1]:I WL[2]:I WL[3]:I WL[4]:I WL[5]:I WL[6]:I WL[7]:I 
*.PININFO WL[8]:I WL[9]:I WL[10]:I WL[11]:I WL[12]:I WL[13]:I WL[14]:I 
*.PININFO WL[15]:I WL[16]:I WL[17]:I WL[18]:I WL[19]:I WL[20]:I WL[21]:I 
*.PININFO WL[22]:I WL[23]:I WL[24]:I WL[25]:I WL[26]:I WL[27]:I WL[28]:I 
*.PININFO WL[29]:I WL[30]:I WL[31]:I WL[32]:I WL[33]:I WL[34]:I WL[35]:I 
*.PININFO WL[36]:I WL[37]:I WL[38]:I WL[39]:I WL[40]:I WL[41]:I WL[42]:I 
*.PININFO WL[43]:I WL[44]:I WL[45]:I WL[46]:I WL[47]:I WL[48]:I WL[49]:I 
*.PININFO WL[50]:I WL[51]:I WL[52]:I WL[53]:I WL[54]:I WL[55]:I WL[56]:I 
*.PININFO WL[57]:I WL[58]:I WL[59]:I WL[60]:I WL[61]:I WL[62]:I WL[63]:I 
*.PININFO WL[64]:I WL[65]:I WL[66]:I WL[67]:I WL[68]:I WL[69]:I WL[70]:I 
*.PININFO WL[71]:I WL[72]:I WL[73]:I WL[74]:I WL[75]:I WL[76]:I WL[77]:I 
*.PININFO WL[78]:I WL[79]:I WL[80]:I WL[81]:I WL[82]:I WL[83]:I WL[84]:I 
*.PININFO WL[85]:I WL[86]:I WL[87]:I WL[88]:I WL[89]:I WL[90]:I WL[91]:I 
*.PININFO WL[92]:I WL[93]:I WL[94]:I WL[95]:I WL[96]:I WL[97]:I WL[98]:I 
*.PININFO WL[99]:I WL[100]:I WL[101]:I WL[102]:I WL[103]:I WL[104]:I WL[105]:I 
*.PININFO WL[106]:I WL[107]:I WL[108]:I WL[109]:I WL[110]:I WL[111]:I 
*.PININFO WL[112]:I WL[113]:I WL[114]:I WL[115]:I WL[116]:I WL[117]:I 
*.PININFO WL[118]:I WL[119]:I WL[120]:I WL[121]:I WL[122]:I WL[123]:I 
*.PININFO WL[124]:I WL[125]:I WL[126]:I WL[127]:I WL[128]:I WL[129]:I 
*.PININFO WL[130]:I WL[131]:I WL[132]:I WL[133]:I WL[134]:I WL[135]:I 
*.PININFO WL[136]:I WL[137]:I WL[138]:I WL[139]:I WL[140]:I WL[141]:I 
*.PININFO WL[142]:I WL[143]:I WL[144]:I WL[145]:I WL[146]:I WL[147]:I 
*.PININFO WL[148]:I WL[149]:I WL[150]:I WL[151]:I WL[152]:I WL[153]:I 
*.PININFO WL[154]:I WL[155]:I WL[156]:I WL[157]:I WL[158]:I WL[159]:I 
*.PININFO WL[160]:I WL[161]:I WL[162]:I WL[163]:I WL[164]:I WL[165]:I 
*.PININFO WL[166]:I WL[167]:I WL[168]:I WL[169]:I WL[170]:I WL[171]:I 
*.PININFO WL[172]:I WL[173]:I WL[174]:I WL[175]:I WL[176]:I WL[177]:I 
*.PININFO WL[178]:I WL[179]:I WL[180]:I WL[181]:I WL[182]:I WL[183]:I 
*.PININFO WL[184]:I WL[185]:I WL[186]:I WL[187]:I WL[188]:I WL[189]:I 
*.PININFO WL[190]:I WL[191]:I WL[192]:I WL[193]:I WL[194]:I WL[195]:I 
*.PININFO WL[196]:I WL[197]:I WL[198]:I WL[199]:I WL[200]:I WL[201]:I 
*.PININFO WL[202]:I WL[203]:I WL[204]:I WL[205]:I WL[206]:I WL[207]:I 
*.PININFO WL[208]:I WL[209]:I WL[210]:I WL[211]:I WL[212]:I WL[213]:I 
*.PININFO WL[214]:I WL[215]:I WL[216]:I WL[217]:I WL[218]:I WL[219]:I 
*.PININFO WL[220]:I WL[221]:I WL[222]:I WL[223]:I WL[224]:I WL[225]:I 
*.PININFO WL[226]:I WL[227]:I WL[228]:I WL[229]:I WL[230]:I WL[231]:I 
*.PININFO WL[232]:I WL[233]:I WL[234]:I WL[235]:I WL[236]:I WL[237]:I 
*.PININFO WL[238]:I WL[239]:I WL[240]:I WL[241]:I WL[242]:I WL[243]:I 
*.PININFO WL[244]:I WL[245]:I WL[246]:I WL[247]:I WL[248]:I WL[249]:I 
*.PININFO WL[250]:I WL[251]:I BL[0]:B BL[1]:B BL[2]:B BL[3]:B BLB[0]:B 
*.PININFO BLB[1]:B BLB[2]:B BLB[3]:B VDDI:B VSSI:B
XMCB_2X4<0> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[0] WL[1] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<1> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[2] WL[3] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<2> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[4] WL[5] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<3> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[6] WL[7] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<4> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[8] WL[9] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<5> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[10] WL[11] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<6> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[12] WL[13] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<7> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[14] WL[15] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<8> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[16] WL[17] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<9> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[18] WL[19] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<10> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[20] WL[21] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<11> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[22] WL[23] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<12> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[24] WL[25] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<13> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[26] WL[27] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<14> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[28] WL[29] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<15> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[30] WL[31] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<16> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[32] WL[33] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<17> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[34] WL[35] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<18> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[36] WL[37] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<19> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[38] WL[39] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<20> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[40] WL[41] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<21> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[42] WL[43] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<22> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[44] WL[45] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<23> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[46] WL[47] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<24> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[48] WL[49] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<25> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[50] WL[51] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<26> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[52] WL[53] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<27> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[54] WL[55] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<28> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[56] WL[57] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<29> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[58] WL[59] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<30> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[60] WL[61] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<31> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[62] WL[63] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<32> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[64] WL[65] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<33> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[66] WL[67] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<34> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[68] WL[69] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<35> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[70] WL[71] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<36> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[72] WL[73] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<37> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[74] WL[75] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<38> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[76] WL[77] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<39> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[78] WL[79] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<40> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[80] WL[81] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<41> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[82] WL[83] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<42> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[84] WL[85] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<43> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[86] WL[87] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<44> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[88] WL[89] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<45> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[90] WL[91] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<46> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[92] WL[93] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<47> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[94] WL[95] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<48> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[96] WL[97] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<49> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[98] WL[99] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<50> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[100] WL[101] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<51> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[102] WL[103] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<52> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[104] WL[105] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<53> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[106] WL[107] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<54> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[108] WL[109] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<55> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[110] WL[111] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<56> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[112] WL[113] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<57> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[114] WL[115] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<58> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[116] WL[117] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<59> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[118] WL[119] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<60> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[120] WL[121] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<61> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[122] WL[123] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<62> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[124] WL[125] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<63> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[126] WL[127] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<64> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[128] WL[129] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<65> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[130] WL[131] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<66> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[132] WL[133] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<67> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[134] WL[135] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<68> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[136] WL[137] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<69> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[138] WL[139] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<70> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[140] WL[141] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<71> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[142] WL[143] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<72> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[144] WL[145] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<73> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[146] WL[147] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<74> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[148] WL[149] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<75> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[150] WL[151] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<76> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[152] WL[153] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<77> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[154] WL[155] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<78> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[156] WL[157] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<79> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[158] WL[159] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<80> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[160] WL[161] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<81> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[162] WL[163] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<82> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[164] WL[165] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<83> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[166] WL[167] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<84> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[168] WL[169] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<85> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[170] WL[171] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<86> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[172] WL[173] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<87> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[174] WL[175] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<88> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[176] WL[177] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<89> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[178] WL[179] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<90> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[180] WL[181] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<91> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[182] WL[183] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<92> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[184] WL[185] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<93> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[186] WL[187] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<94> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[188] WL[189] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<95> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[190] WL[191] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<96> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[192] WL[193] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<97> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[194] WL[195] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<98> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[196] WL[197] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<99> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[198] WL[199] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<100> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[200] WL[201] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<101> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[202] WL[203] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<102> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[204] WL[205] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<103> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[206] WL[207] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<104> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[208] WL[209] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<105> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[210] WL[211] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<106> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[212] WL[213] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<107> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[214] WL[215] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<108> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[216] WL[217] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<109> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[218] WL[219] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<110> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[220] WL[221] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<111> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[222] WL[223] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<112> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[224] WL[225] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<113> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[226] WL[227] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<114> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[228] WL[229] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<115> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[230] WL[231] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<116> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[232] WL[233] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<117> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[234] WL[235] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<118> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[236] WL[237] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<119> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[238] WL[239] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<120> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[240] WL[241] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<121> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[242] WL[243] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<122> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[244] WL[245] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<123> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[246] WL[247] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<124> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[248] WL[249] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<125> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[250] WL[251] S1AHSF400W40_MCB_2X4_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    MCB_124X4_SB_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_124X4_SB_CHAR BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] 
+ VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] 
+ WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] 
+ WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] 
+ WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] 
+ WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] 
+ WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] WL[64] WL[65] 
+ WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] 
+ WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] 
+ WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] 
+ WL[99] WL[100] WL[101] WL[102] WL[103] WL[104] WL[105] WL[106] WL[107] 
+ WL[108] WL[109] WL[110] WL[111] WL[112] WL[113] WL[114] WL[115] WL[116] 
+ WL[117] WL[118] WL[119] WL[120] WL[121] WL[122] WL[123]
*.PININFO WL[0]:I WL[1]:I WL[2]:I WL[3]:I WL[4]:I WL[5]:I WL[6]:I WL[7]:I 
*.PININFO WL[8]:I WL[9]:I WL[10]:I WL[11]:I WL[12]:I WL[13]:I WL[14]:I 
*.PININFO WL[15]:I WL[16]:I WL[17]:I WL[18]:I WL[19]:I WL[20]:I WL[21]:I 
*.PININFO WL[22]:I WL[23]:I WL[24]:I WL[25]:I WL[26]:I WL[27]:I WL[28]:I 
*.PININFO WL[29]:I WL[30]:I WL[31]:I WL[32]:I WL[33]:I WL[34]:I WL[35]:I 
*.PININFO WL[36]:I WL[37]:I WL[38]:I WL[39]:I WL[40]:I WL[41]:I WL[42]:I 
*.PININFO WL[43]:I WL[44]:I WL[45]:I WL[46]:I WL[47]:I WL[48]:I WL[49]:I 
*.PININFO WL[50]:I WL[51]:I WL[52]:I WL[53]:I WL[54]:I WL[55]:I WL[56]:I 
*.PININFO WL[57]:I WL[58]:I WL[59]:I WL[60]:I WL[61]:I WL[62]:I WL[63]:I 
*.PININFO WL[64]:I WL[65]:I WL[66]:I WL[67]:I WL[68]:I WL[69]:I WL[70]:I 
*.PININFO WL[71]:I WL[72]:I WL[73]:I WL[74]:I WL[75]:I WL[76]:I WL[77]:I 
*.PININFO WL[78]:I WL[79]:I WL[80]:I WL[81]:I WL[82]:I WL[83]:I WL[84]:I 
*.PININFO WL[85]:I WL[86]:I WL[87]:I WL[88]:I WL[89]:I WL[90]:I WL[91]:I 
*.PININFO WL[92]:I WL[93]:I WL[94]:I WL[95]:I WL[96]:I WL[97]:I WL[98]:I 
*.PININFO WL[99]:I WL[100]:I WL[101]:I WL[102]:I WL[103]:I WL[104]:I WL[105]:I 
*.PININFO WL[106]:I WL[107]:I WL[108]:I WL[109]:I WL[110]:I WL[111]:I 
*.PININFO WL[112]:I WL[113]:I WL[114]:I WL[115]:I WL[116]:I WL[117]:I 
*.PININFO WL[118]:I WL[119]:I WL[120]:I WL[121]:I WL[122]:I WL[123]:I BL[0]:B 
*.PININFO BL[1]:B BL[2]:B BL[3]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B VDDI:B 
*.PININFO VSSI:B
XMCB_2X4<0> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[0] WL[1] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<1> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[2] WL[3] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<2> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[4] WL[5] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<3> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[6] WL[7] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<4> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[8] WL[9] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<5> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[10] WL[11] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<6> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[12] WL[13] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<7> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[14] WL[15] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<8> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[16] WL[17] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<9> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[18] WL[19] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<10> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[20] WL[21] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<11> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[22] WL[23] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<12> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[24] WL[25] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<13> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[26] WL[27] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<14> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[28] WL[29] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<15> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[30] WL[31] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<16> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[32] WL[33] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<17> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[34] WL[35] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<18> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[36] WL[37] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<19> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[38] WL[39] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<20> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[40] WL[41] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<21> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[42] WL[43] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<22> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[44] WL[45] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<23> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[46] WL[47] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<24> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[48] WL[49] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<25> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[50] WL[51] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<26> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[52] WL[53] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<27> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[54] WL[55] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<28> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[56] WL[57] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<29> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[58] WL[59] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<30> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[60] WL[61] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<31> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[62] WL[63] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<32> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[64] WL[65] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<33> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[66] WL[67] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<34> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[68] WL[69] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<35> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[70] WL[71] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<36> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[72] WL[73] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<37> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[74] WL[75] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<38> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[76] WL[77] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<39> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[78] WL[79] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<40> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[80] WL[81] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<41> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[82] WL[83] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<42> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[84] WL[85] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<43> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[86] WL[87] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<44> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[88] WL[89] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<45> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[90] WL[91] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<46> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[92] WL[93] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<47> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[94] WL[95] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<48> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[96] WL[97] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<49> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[98] WL[99] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<50> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[100] WL[101] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<51> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[102] WL[103] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<52> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[104] WL[105] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<53> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[106] WL[107] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<54> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[108] WL[109] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<55> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[110] WL[111] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<56> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[112] WL[113] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<57> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[114] WL[115] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<58> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[116] WL[117] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<59> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[118] WL[119] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<60> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[120] WL[121] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<61> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[122] WL[123] S1AHSF400W40_MCB_2X4_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    MCB_12X4_SB_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_12X4_SB_CHAR BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] 
+ VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] 
+ WL[11]
*.PININFO WL[0]:I WL[1]:I WL[2]:I WL[3]:I WL[4]:I WL[5]:I WL[6]:I WL[7]:I 
*.PININFO WL[8]:I WL[9]:I WL[10]:I WL[11]:I BL[0]:B BL[1]:B BL[2]:B BL[3]:B 
*.PININFO BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B VDDI:B VSSI:B
XMCB_2X4<0> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[0] WL[1] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<1> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[2] WL[3] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<2> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[4] WL[5] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<3> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[6] WL[7] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<4> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[8] WL[9] S1AHSF400W40_MCB_2X4_SB
XMCB_2X4<5> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] VDDI VSSI 
+ WL[10] WL[11] S1AHSF400W40_MCB_2X4_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_ARR_BLLD_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_ARR_BLLD_SIM BLB_BT[0] BLB_TP[0] BL_BT[0] BL_TP[0] VDDI VSSI
*.PININFO BLB_BT[0]:B BLB_TP[0]:B BL_BT[0]:B BL_TP[0]:B VDDI:B VSSI:B
XI43 NET062[0] NET062[1] NET062[2] NET062[3] NET049[0] NET049[1] NET049[2] 
+ NET049[3] NET054 NET061 NET070[0] NET070[1] NET070[2] NET070[3] NET070[4] 
+ NET070[5] NET070[6] NET070[7] NET070[8] NET070[9] NET070[10] NET070[11] 
+ NET070[12] NET070[13] NET070[14] NET070[15] NET070[16] NET070[17] NET070[18] 
+ NET070[19] NET070[20] NET070[21] NET070[22] NET070[23] NET070[24] NET070[25] 
+ NET070[26] NET070[27] NET070[28] NET070[29] NET070[30] NET070[31] NET070[32] 
+ NET070[33] NET070[34] NET070[35] NET070[36] NET070[37] NET070[38] NET070[39] 
+ NET070[40] NET070[41] NET070[42] NET070[43] NET070[44] NET070[45] NET070[46] 
+ NET070[47] NET070[48] NET070[49] NET070[50] NET070[51] NET070[52] NET070[53] 
+ NET070[54] NET070[55] NET070[56] NET070[57] NET070[58] NET070[59] NET070[60] 
+ NET070[61] S1AHSF400W40_MCB_62X4_SB_CHAR
XI42 NET042[0] NET042[1] NET042[2] NET042[3] NET02[0] NET02[1] NET02[2] 
+ NET02[3] NET060 NET038 NET075[0] NET075[1] NET075[2] NET075[3] NET075[4] 
+ NET075[5] NET075[6] NET075[7] NET075[8] NET075[9] NET075[10] NET075[11] 
+ NET075[12] NET075[13] NET075[14] NET075[15] NET075[16] NET075[17] NET075[18] 
+ NET075[19] NET075[20] NET075[21] NET075[22] NET075[23] NET075[24] NET075[25] 
+ NET075[26] NET075[27] NET075[28] NET075[29] NET075[30] NET075[31] NET075[32] 
+ NET075[33] NET075[34] NET075[35] NET075[36] NET075[37] NET075[38] NET075[39] 
+ NET075[40] NET075[41] NET075[42] NET075[43] NET075[44] NET075[45] NET075[46] 
+ NET075[47] NET075[48] NET075[49] NET075[50] NET075[51] NET075[52] NET075[53] 
+ NET075[54] NET075[55] NET075[56] NET075[57] NET075[58] NET075[59] 
+ S1AHSF400W40_MCB_60X4_SB_CHAR
XI44 NET056[0] NET056[1] NET056[2] NET056[3] NET057[0] NET057[1] NET057[2] 
+ NET057[3] NET055 NET059 NET080[0] NET080[1] NET080[2] NET080[3] NET080[4] 
+ NET080[5] NET080[6] NET080[7] NET080[8] NET080[9] NET080[10] NET080[11] 
+ NET080[12] NET080[13] NET080[14] NET080[15] NET080[16] NET080[17] NET080[18] 
+ NET080[19] NET080[20] NET080[21] NET080[22] NET080[23] NET080[24] NET080[25] 
+ NET080[26] NET080[27] NET080[28] NET080[29] NET080[30] NET080[31] NET080[32] 
+ NET080[33] NET080[34] NET080[35] NET080[36] NET080[37] NET080[38] NET080[39] 
+ NET080[40] NET080[41] NET080[42] NET080[43] NET080[44] NET080[45] NET080[46] 
+ NET080[47] NET080[48] NET080[49] NET080[50] NET080[51] NET080[52] NET080[53] 
+ NET080[54] NET080[55] NET080[56] NET080[57] NET080[58] NET080[59] NET080[60] 
+ NET080[61] NET080[62] NET080[63] NET080[64] NET080[65] NET080[66] NET080[67] 
+ NET080[68] NET080[69] NET080[70] NET080[71] NET080[72] NET080[73] NET080[74] 
+ NET080[75] NET080[76] NET080[77] NET080[78] NET080[79] NET080[80] NET080[81] 
+ NET080[82] NET080[83] NET080[84] NET080[85] NET080[86] NET080[87] NET080[88] 
+ NET080[89] NET080[90] NET080[91] NET080[92] NET080[93] NET080[94] NET080[95] 
+ NET080[96] NET080[97] NET080[98] NET080[99] NET080[100] NET080[101] 
+ NET080[102] NET080[103] NET080[104] NET080[105] NET080[106] NET080[107] 
+ NET080[108] NET080[109] NET080[110] NET080[111] NET080[112] NET080[113] 
+ NET080[114] NET080[115] NET080[116] NET080[117] NET080[118] NET080[119] 
+ NET080[120] NET080[121] NET080[122] NET080[123] NET080[124] NET080[125] 
+ NET080[126] NET080[127] NET080[128] NET080[129] NET080[130] NET080[131] 
+ NET080[132] NET080[133] NET080[134] NET080[135] NET080[136] NET080[137] 
+ NET080[138] NET080[139] NET080[140] NET080[141] NET080[142] NET080[143] 
+ NET080[144] NET080[145] NET080[146] NET080[147] NET080[148] NET080[149] 
+ NET080[150] NET080[151] NET080[152] NET080[153] NET080[154] NET080[155] 
+ NET080[156] NET080[157] NET080[158] NET080[159] NET080[160] NET080[161] 
+ NET080[162] NET080[163] NET080[164] NET080[165] NET080[166] NET080[167] 
+ NET080[168] NET080[169] NET080[170] NET080[171] NET080[172] NET080[173] 
+ NET080[174] NET080[175] NET080[176] NET080[177] NET080[178] NET080[179] 
+ NET080[180] NET080[181] NET080[182] NET080[183] NET080[184] NET080[185] 
+ NET080[186] NET080[187] NET080[188] NET080[189] NET080[190] NET080[191] 
+ NET080[192] NET080[193] NET080[194] NET080[195] NET080[196] NET080[197] 
+ NET080[198] NET080[199] NET080[200] NET080[201] NET080[202] NET080[203] 
+ NET080[204] NET080[205] NET080[206] NET080[207] NET080[208] NET080[209] 
+ NET080[210] NET080[211] NET080[212] NET080[213] NET080[214] NET080[215] 
+ NET080[216] NET080[217] NET080[218] NET080[219] NET080[220] NET080[221] 
+ NET080[222] NET080[223] NET080[224] NET080[225] NET080[226] NET080[227] 
+ NET080[228] NET080[229] NET080[230] NET080[231] NET080[232] NET080[233] 
+ NET080[234] NET080[235] NET080[236] NET080[237] NET080[238] NET080[239] 
+ NET080[240] NET080[241] NET080[242] NET080[243] NET080[244] NET080[245] 
+ NET080[246] NET080[247] NET080[248] NET080[249] NET080[250] NET080[251] 
+ NET080[252] NET080[253] NET080[254] NET080[255] NET080[256] NET080[257] 
+ NET080[258] NET080[259] NET080[260] NET080[261] NET080[262] NET080[263] 
+ NET080[264] NET080[265] NET080[266] NET080[267] NET080[268] NET080[269] 
+ NET080[270] NET080[271] NET080[272] NET080[273] NET080[274] NET080[275] 
+ NET080[276] NET080[277] NET080[278] NET080[279] NET080[280] NET080[281] 
+ NET080[282] NET080[283] NET080[284] NET080[285] NET080[286] NET080[287] 
+ NET080[288] NET080[289] NET080[290] NET080[291] NET080[292] NET080[293] 
+ NET080[294] NET080[295] NET080[296] NET080[297] NET080[298] NET080[299] 
+ NET080[300] NET080[301] NET080[302] NET080[303] NET080[304] NET080[305] 
+ NET080[306] NET080[307] NET080[308] NET080[309] NET080[310] NET080[311] 
+ NET080[312] NET080[313] NET080[314] NET080[315] NET080[316] NET080[317] 
+ NET080[318] NET080[319] NET080[320] NET080[321] NET080[322] NET080[323] 
+ NET080[324] NET080[325] NET080[326] NET080[327] NET080[328] NET080[329] 
+ NET080[330] NET080[331] NET080[332] NET080[333] NET080[334] NET080[335] 
+ NET080[336] NET080[337] NET080[338] NET080[339] NET080[340] NET080[341] 
+ NET080[342] NET080[343] NET080[344] NET080[345] NET080[346] NET080[347] 
+ NET080[348] NET080[349] NET080[350] NET080[351] NET080[352] NET080[353] 
+ NET080[354] NET080[355] NET080[356] NET080[357] NET080[358] NET080[359] 
+ NET080[360] NET080[361] NET080[362] NET080[363] NET080[364] NET080[365] 
+ NET080[366] NET080[367] NET080[368] NET080[369] NET080[370] NET080[371] 
+ NET080[372] NET080[373] NET080[374] NET080[375] NET080[376] NET080[377] 
+ NET080[378] NET080[379] S1AHSF400W40_MCB_380X4_SB_CHAR
XI45 NET024[0] NET024[1] NET024[2] NET024[3] NET023[0] NET023[1] NET023[2] 
+ NET023[3] NET046 NET063 NET085[0] NET085[1] NET085[2] NET085[3] NET085[4] 
+ NET085[5] NET085[6] NET085[7] NET085[8] NET085[9] NET085[10] NET085[11] 
+ NET085[12] NET085[13] NET085[14] NET085[15] NET085[16] NET085[17] NET085[18] 
+ NET085[19] NET085[20] NET085[21] NET085[22] NET085[23] NET085[24] NET085[25] 
+ NET085[26] NET085[27] NET085[28] NET085[29] NET085[30] NET085[31] NET085[32] 
+ NET085[33] NET085[34] NET085[35] NET085[36] NET085[37] NET085[38] NET085[39] 
+ NET085[40] NET085[41] NET085[42] NET085[43] NET085[44] NET085[45] NET085[46] 
+ NET085[47] NET085[48] NET085[49] NET085[50] NET085[51] NET085[52] NET085[53] 
+ NET085[54] NET085[55] NET085[56] NET085[57] NET085[58] NET085[59] NET085[60] 
+ NET085[61] NET085[62] NET085[63] NET085[64] NET085[65] NET085[66] NET085[67] 
+ NET085[68] NET085[69] NET085[70] NET085[71] NET085[72] NET085[73] NET085[74] 
+ NET085[75] NET085[76] NET085[77] NET085[78] NET085[79] NET085[80] NET085[81] 
+ NET085[82] NET085[83] NET085[84] NET085[85] NET085[86] NET085[87] NET085[88] 
+ NET085[89] NET085[90] NET085[91] NET085[92] NET085[93] NET085[94] NET085[95] 
+ NET085[96] NET085[97] NET085[98] NET085[99] NET085[100] NET085[101] 
+ NET085[102] NET085[103] NET085[104] NET085[105] NET085[106] NET085[107] 
+ NET085[108] NET085[109] NET085[110] NET085[111] NET085[112] NET085[113] 
+ NET085[114] NET085[115] NET085[116] NET085[117] NET085[118] NET085[119] 
+ NET085[120] NET085[121] NET085[122] NET085[123] NET085[124] NET085[125] 
+ NET085[126] NET085[127] NET085[128] NET085[129] NET085[130] NET085[131] 
+ NET085[132] NET085[133] NET085[134] NET085[135] NET085[136] NET085[137] 
+ NET085[138] NET085[139] NET085[140] NET085[141] NET085[142] NET085[143] 
+ NET085[144] NET085[145] NET085[146] NET085[147] NET085[148] NET085[149] 
+ NET085[150] NET085[151] NET085[152] NET085[153] NET085[154] NET085[155] 
+ NET085[156] NET085[157] NET085[158] NET085[159] NET085[160] NET085[161] 
+ NET085[162] NET085[163] NET085[164] NET085[165] NET085[166] NET085[167] 
+ NET085[168] NET085[169] NET085[170] NET085[171] NET085[172] NET085[173] 
+ NET085[174] NET085[175] NET085[176] NET085[177] NET085[178] NET085[179] 
+ NET085[180] NET085[181] NET085[182] NET085[183] NET085[184] NET085[185] 
+ NET085[186] NET085[187] NET085[188] NET085[189] NET085[190] NET085[191] 
+ NET085[192] NET085[193] NET085[194] NET085[195] NET085[196] NET085[197] 
+ NET085[198] NET085[199] NET085[200] NET085[201] NET085[202] NET085[203] 
+ NET085[204] NET085[205] NET085[206] NET085[207] NET085[208] NET085[209] 
+ NET085[210] NET085[211] NET085[212] NET085[213] NET085[214] NET085[215] 
+ NET085[216] NET085[217] NET085[218] NET085[219] NET085[220] NET085[221] 
+ NET085[222] NET085[223] NET085[224] NET085[225] NET085[226] NET085[227] 
+ NET085[228] NET085[229] NET085[230] NET085[231] NET085[232] NET085[233] 
+ NET085[234] NET085[235] NET085[236] NET085[237] NET085[238] NET085[239] 
+ NET085[240] NET085[241] NET085[242] NET085[243] NET085[244] NET085[245] 
+ NET085[246] NET085[247] NET085[248] NET085[249] NET085[250] NET085[251] 
+ NET085[252] NET085[253] NET085[254] NET085[255] NET085[256] NET085[257] 
+ NET085[258] NET085[259] NET085[260] NET085[261] NET085[262] NET085[263] 
+ NET085[264] NET085[265] NET085[266] NET085[267] NET085[268] NET085[269] 
+ NET085[270] NET085[271] NET085[272] NET085[273] NET085[274] NET085[275] 
+ NET085[276] NET085[277] NET085[278] NET085[279] NET085[280] NET085[281] 
+ NET085[282] NET085[283] NET085[284] NET085[285] NET085[286] NET085[287] 
+ NET085[288] NET085[289] NET085[290] NET085[291] NET085[292] NET085[293] 
+ NET085[294] NET085[295] NET085[296] NET085[297] NET085[298] NET085[299] 
+ NET085[300] NET085[301] NET085[302] NET085[303] NET085[304] NET085[305] 
+ NET085[306] NET085[307] NET085[308] NET085[309] NET085[310] NET085[311] 
+ NET085[312] NET085[313] NET085[314] NET085[315] NET085[316] NET085[317] 
+ NET085[318] NET085[319] NET085[320] NET085[321] NET085[322] NET085[323] 
+ NET085[324] NET085[325] NET085[326] NET085[327] NET085[328] NET085[329] 
+ NET085[330] NET085[331] NET085[332] NET085[333] NET085[334] NET085[335] 
+ NET085[336] NET085[337] NET085[338] NET085[339] NET085[340] NET085[341] 
+ NET085[342] NET085[343] NET085[344] NET085[345] NET085[346] NET085[347] 
+ NET085[348] NET085[349] NET085[350] NET085[351] NET085[352] NET085[353] 
+ NET085[354] NET085[355] NET085[356] NET085[357] NET085[358] NET085[359] 
+ NET085[360] NET085[361] NET085[362] NET085[363] NET085[364] NET085[365] 
+ NET085[366] NET085[367] NET085[368] NET085[369] NET085[370] NET085[371] 
+ NET085[372] NET085[373] NET085[374] NET085[375] NET085[376] NET085[377] 
+ NET085[378] NET085[379] NET085[380] NET085[381] S1AHSF400W40_MCB_382X4_SB_CHAR
XI39 NET019[0] NET019[1] NET019[2] NET019[3] NET018[0] NET018[1] NET018[2] 
+ NET018[3] NET020 NET021 NET032[0] NET032[1] NET032[2] NET032[3] NET032[4] 
+ NET032[5] NET032[6] NET032[7] NET032[8] NET032[9] NET032[10] NET032[11] 
+ NET032[12] NET032[13] NET032[14] NET032[15] NET032[16] NET032[17] NET032[18] 
+ NET032[19] NET032[20] NET032[21] NET032[22] NET032[23] NET032[24] NET032[25] 
+ NET032[26] NET032[27] NET032[28] NET032[29] NET032[30] NET032[31] NET032[32] 
+ NET032[33] NET032[34] NET032[35] NET032[36] NET032[37] NET032[38] NET032[39] 
+ NET032[40] NET032[41] NET032[42] NET032[43] NET032[44] NET032[45] NET032[46] 
+ NET032[47] NET032[48] NET032[49] NET032[50] NET032[51] NET032[52] NET032[53] 
+ NET032[54] NET032[55] NET032[56] NET032[57] NET032[58] NET032[59] NET032[60] 
+ NET032[61] NET032[62] NET032[63] NET032[64] NET032[65] NET032[66] NET032[67] 
+ NET032[68] NET032[69] NET032[70] NET032[71] NET032[72] NET032[73] NET032[74] 
+ NET032[75] NET032[76] NET032[77] NET032[78] NET032[79] NET032[80] NET032[81] 
+ NET032[82] NET032[83] NET032[84] NET032[85] NET032[86] NET032[87] NET032[88] 
+ NET032[89] NET032[90] NET032[91] NET032[92] NET032[93] NET032[94] NET032[95] 
+ NET032[96] NET032[97] NET032[98] NET032[99] NET032[100] NET032[101] 
+ NET032[102] NET032[103] NET032[104] NET032[105] NET032[106] NET032[107] 
+ NET032[108] NET032[109] NET032[110] NET032[111] NET032[112] NET032[113] 
+ NET032[114] NET032[115] NET032[116] NET032[117] NET032[118] NET032[119] 
+ NET032[120] NET032[121] NET032[122] NET032[123] NET032[124] NET032[125] 
+ NET032[126] NET032[127] NET032[128] NET032[129] NET032[130] NET032[131] 
+ NET032[132] NET032[133] NET032[134] NET032[135] NET032[136] NET032[137] 
+ NET032[138] NET032[139] NET032[140] NET032[141] NET032[142] NET032[143] 
+ NET032[144] NET032[145] NET032[146] NET032[147] NET032[148] NET032[149] 
+ NET032[150] NET032[151] NET032[152] NET032[153] NET032[154] NET032[155] 
+ NET032[156] NET032[157] NET032[158] NET032[159] NET032[160] NET032[161] 
+ NET032[162] NET032[163] NET032[164] NET032[165] NET032[166] NET032[167] 
+ NET032[168] NET032[169] NET032[170] NET032[171] NET032[172] NET032[173] 
+ NET032[174] NET032[175] NET032[176] NET032[177] NET032[178] NET032[179] 
+ NET032[180] NET032[181] NET032[182] NET032[183] NET032[184] NET032[185] 
+ NET032[186] NET032[187] NET032[188] NET032[189] NET032[190] NET032[191] 
+ NET032[192] NET032[193] NET032[194] NET032[195] NET032[196] NET032[197] 
+ NET032[198] NET032[199] NET032[200] NET032[201] NET032[202] NET032[203] 
+ NET032[204] NET032[205] NET032[206] NET032[207] NET032[208] NET032[209] 
+ NET032[210] NET032[211] NET032[212] NET032[213] NET032[214] NET032[215] 
+ NET032[216] NET032[217] NET032[218] NET032[219] NET032[220] NET032[221] 
+ NET032[222] NET032[223] NET032[224] NET032[225] NET032[226] NET032[227] 
+ NET032[228] NET032[229] NET032[230] NET032[231] NET032[232] NET032[233] 
+ NET032[234] NET032[235] NET032[236] NET032[237] NET032[238] NET032[239] 
+ NET032[240] NET032[241] NET032[242] NET032[243] NET032[244] NET032[245] 
+ NET032[246] NET032[247] NET032[248] NET032[249] NET032[250] NET032[251] 
+ NET032[252] NET032[253] NET032[254] NET032[255] NET032[256] NET032[257] 
+ NET032[258] NET032[259] NET032[260] NET032[261] NET032[262] NET032[263] 
+ NET032[264] NET032[265] NET032[266] NET032[267] NET032[268] NET032[269] 
+ NET032[270] NET032[271] NET032[272] NET032[273] NET032[274] NET032[275] 
+ NET032[276] NET032[277] NET032[278] NET032[279] NET032[280] NET032[281] 
+ NET032[282] NET032[283] NET032[284] NET032[285] NET032[286] NET032[287] 
+ NET032[288] NET032[289] NET032[290] NET032[291] NET032[292] NET032[293] 
+ NET032[294] NET032[295] NET032[296] NET032[297] NET032[298] NET032[299] 
+ NET032[300] NET032[301] NET032[302] NET032[303] NET032[304] NET032[305] 
+ NET032[306] NET032[307] NET032[308] NET032[309] NET032[310] NET032[311] 
+ NET032[312] NET032[313] NET032[314] NET032[315] NET032[316] NET032[317] 
+ NET032[318] NET032[319] NET032[320] NET032[321] NET032[322] NET032[323] 
+ NET032[324] NET032[325] NET032[326] NET032[327] NET032[328] NET032[329] 
+ NET032[330] NET032[331] NET032[332] NET032[333] NET032[334] NET032[335] 
+ NET032[336] NET032[337] NET032[338] NET032[339] NET032[340] NET032[341] 
+ NET032[342] NET032[343] NET032[344] NET032[345] NET032[346] NET032[347] 
+ NET032[348] NET032[349] NET032[350] NET032[351] NET032[352] NET032[353] 
+ NET032[354] NET032[355] NET032[356] NET032[357] NET032[358] NET032[359] 
+ NET032[360] NET032[361] NET032[362] NET032[363] NET032[364] NET032[365] 
+ NET032[366] NET032[367] NET032[368] NET032[369] NET032[370] NET032[371] 
+ NET032[372] NET032[373] NET032[374] NET032[375] NET032[376] NET032[377] 
+ NET032[378] NET032[379] NET032[380] NET032[381] NET032[382] NET032[383] 
+ NET032[384] NET032[385] NET032[386] NET032[387] NET032[388] NET032[389] 
+ NET032[390] NET032[391] NET032[392] NET032[393] NET032[394] NET032[395] 
+ NET032[396] NET032[397] NET032[398] NET032[399] NET032[400] NET032[401] 
+ NET032[402] NET032[403] NET032[404] NET032[405] NET032[406] NET032[407] 
+ NET032[408] NET032[409] NET032[410] NET032[411] NET032[412] NET032[413] 
+ NET032[414] NET032[415] NET032[416] NET032[417] NET032[418] NET032[419] 
+ NET032[420] NET032[421] NET032[422] NET032[423] NET032[424] NET032[425] 
+ NET032[426] NET032[427] NET032[428] NET032[429] NET032[430] NET032[431] 
+ NET032[432] NET032[433] NET032[434] NET032[435] NET032[436] NET032[437] 
+ NET032[438] NET032[439] NET032[440] NET032[441] NET032[442] NET032[443] 
+ NET032[444] NET032[445] NET032[446] NET032[447] NET032[448] NET032[449] 
+ NET032[450] NET032[451] NET032[452] NET032[453] NET032[454] NET032[455] 
+ NET032[456] NET032[457] NET032[458] NET032[459] NET032[460] NET032[461] 
+ NET032[462] NET032[463] NET032[464] NET032[465] NET032[466] NET032[467] 
+ NET032[468] NET032[469] NET032[470] NET032[471] NET032[472] NET032[473] 
+ NET032[474] NET032[475] NET032[476] NET032[477] NET032[478] NET032[479] 
+ NET032[480] NET032[481] NET032[482] NET032[483] NET032[484] NET032[485] 
+ NET032[486] NET032[487] NET032[488] NET032[489] NET032[490] NET032[491] 
+ NET032[492] NET032[493] NET032[494] NET032[495] NET032[496] NET032[497] 
+ NET032[498] NET032[499] NET032[500] NET032[501] NET032[502] NET032[503] 
+ NET032[504] NET032[505] NET032[506] NET032[507] S1AHSF400W40_MCB_508X4_SB_CHAR
XI41 NET029[0] NET029[1] NET029[2] NET029[3] NET026[0] NET026[1] NET026[2] 
+ NET026[3] NET027 NET03 NET025[0] NET025[1] NET025[2] NET025[3] NET025[4] 
+ NET025[5] NET025[6] NET025[7] NET025[8] NET025[9] NET025[10] NET025[11] 
+ NET025[12] NET025[13] NET025[14] NET025[15] NET025[16] NET025[17] NET025[18] 
+ NET025[19] NET025[20] NET025[21] NET025[22] NET025[23] NET025[24] NET025[25] 
+ NET025[26] NET025[27] NET025[28] NET025[29] NET025[30] NET025[31] NET025[32] 
+ NET025[33] NET025[34] NET025[35] NET025[36] NET025[37] NET025[38] NET025[39] 
+ NET025[40] NET025[41] NET025[42] NET025[43] NET025[44] NET025[45] NET025[46] 
+ NET025[47] NET025[48] NET025[49] NET025[50] NET025[51] NET025[52] NET025[53] 
+ NET025[54] NET025[55] NET025[56] NET025[57] NET025[58] NET025[59] NET025[60] 
+ NET025[61] NET025[62] NET025[63] NET025[64] NET025[65] NET025[66] NET025[67] 
+ NET025[68] NET025[69] NET025[70] NET025[71] NET025[72] NET025[73] NET025[74] 
+ NET025[75] NET025[76] NET025[77] NET025[78] NET025[79] NET025[80] NET025[81] 
+ NET025[82] NET025[83] NET025[84] NET025[85] NET025[86] NET025[87] NET025[88] 
+ NET025[89] NET025[90] NET025[91] NET025[92] NET025[93] NET025[94] NET025[95] 
+ NET025[96] NET025[97] NET025[98] NET025[99] NET025[100] NET025[101] 
+ NET025[102] NET025[103] NET025[104] NET025[105] NET025[106] NET025[107] 
+ NET025[108] NET025[109] NET025[110] NET025[111] NET025[112] NET025[113] 
+ NET025[114] NET025[115] NET025[116] NET025[117] NET025[118] NET025[119] 
+ NET025[120] NET025[121] NET025[122] NET025[123] NET025[124] NET025[125] 
+ NET025[126] NET025[127] NET025[128] NET025[129] NET025[130] NET025[131] 
+ NET025[132] NET025[133] NET025[134] NET025[135] NET025[136] NET025[137] 
+ NET025[138] NET025[139] NET025[140] NET025[141] NET025[142] NET025[143] 
+ NET025[144] NET025[145] NET025[146] NET025[147] NET025[148] NET025[149] 
+ NET025[150] NET025[151] NET025[152] NET025[153] NET025[154] NET025[155] 
+ NET025[156] NET025[157] NET025[158] NET025[159] NET025[160] NET025[161] 
+ NET025[162] NET025[163] NET025[164] NET025[165] NET025[166] NET025[167] 
+ NET025[168] NET025[169] NET025[170] NET025[171] NET025[172] NET025[173] 
+ NET025[174] NET025[175] NET025[176] NET025[177] NET025[178] NET025[179] 
+ NET025[180] NET025[181] NET025[182] NET025[183] NET025[184] NET025[185] 
+ NET025[186] NET025[187] NET025[188] NET025[189] NET025[190] NET025[191] 
+ NET025[192] NET025[193] NET025[194] NET025[195] NET025[196] NET025[197] 
+ NET025[198] NET025[199] NET025[200] NET025[201] NET025[202] NET025[203] 
+ NET025[204] NET025[205] NET025[206] NET025[207] NET025[208] NET025[209] 
+ NET025[210] NET025[211] NET025[212] NET025[213] NET025[214] NET025[215] 
+ NET025[216] NET025[217] NET025[218] NET025[219] NET025[220] NET025[221] 
+ NET025[222] NET025[223] NET025[224] NET025[225] NET025[226] NET025[227] 
+ NET025[228] NET025[229] NET025[230] NET025[231] NET025[232] NET025[233] 
+ NET025[234] NET025[235] NET025[236] NET025[237] NET025[238] NET025[239] 
+ NET025[240] NET025[241] NET025[242] NET025[243] NET025[244] NET025[245] 
+ NET025[246] NET025[247] NET025[248] NET025[249] NET025[250] NET025[251] 
+ NET025[252] NET025[253] S1AHSF400W40_MCB_254X4_SB_CHAR
XI40 NET06[0] NET06[1] NET06[2] NET06[3] NET01[0] NET01[1] NET01[2] NET01[3] 
+ NET04 NET05 NET022[0] NET022[1] NET022[2] NET022[3] NET022[4] NET022[5] 
+ NET022[6] NET022[7] NET022[8] NET022[9] NET022[10] NET022[11] NET022[12] 
+ NET022[13] NET022[14] NET022[15] NET022[16] NET022[17] NET022[18] NET022[19] 
+ NET022[20] NET022[21] NET022[22] NET022[23] NET022[24] NET022[25] NET022[26] 
+ NET022[27] NET022[28] NET022[29] NET022[30] NET022[31] NET022[32] NET022[33] 
+ NET022[34] NET022[35] NET022[36] NET022[37] NET022[38] NET022[39] NET022[40] 
+ NET022[41] NET022[42] NET022[43] NET022[44] NET022[45] NET022[46] NET022[47] 
+ NET022[48] NET022[49] NET022[50] NET022[51] NET022[52] NET022[53] NET022[54] 
+ NET022[55] NET022[56] NET022[57] NET022[58] NET022[59] NET022[60] NET022[61] 
+ NET022[62] NET022[63] NET022[64] NET022[65] NET022[66] NET022[67] NET022[68] 
+ NET022[69] NET022[70] NET022[71] NET022[72] NET022[73] NET022[74] NET022[75] 
+ NET022[76] NET022[77] NET022[78] NET022[79] NET022[80] NET022[81] NET022[82] 
+ NET022[83] NET022[84] NET022[85] NET022[86] NET022[87] NET022[88] NET022[89] 
+ NET022[90] NET022[91] NET022[92] NET022[93] NET022[94] NET022[95] NET022[96] 
+ NET022[97] NET022[98] NET022[99] NET022[100] NET022[101] NET022[102] 
+ NET022[103] NET022[104] NET022[105] NET022[106] NET022[107] NET022[108] 
+ NET022[109] NET022[110] NET022[111] NET022[112] NET022[113] NET022[114] 
+ NET022[115] NET022[116] NET022[117] NET022[118] NET022[119] NET022[120] 
+ NET022[121] NET022[122] NET022[123] NET022[124] NET022[125] 
+ S1AHSF400W40_MCB_126X4_SB_CHAR
XI38 NET09[0] NET09[1] NET09[2] NET09[3] NET08[0] NET08[1] NET08[2] NET08[3] 
+ NET010 NET011 NET017[0] NET017[1] NET017[2] NET017[3] NET017[4] NET017[5] 
+ NET017[6] NET017[7] NET017[8] NET017[9] NET017[10] NET017[11] NET017[12] 
+ NET017[13] NET017[14] NET017[15] NET017[16] NET017[17] NET017[18] NET017[19] 
+ NET017[20] NET017[21] NET017[22] NET017[23] NET017[24] NET017[25] NET017[26] 
+ NET017[27] NET017[28] NET017[29] NET017[30] NET017[31] NET017[32] NET017[33] 
+ NET017[34] NET017[35] NET017[36] NET017[37] NET017[38] NET017[39] NET017[40] 
+ NET017[41] NET017[42] NET017[43] NET017[44] NET017[45] NET017[46] NET017[47] 
+ NET017[48] NET017[49] NET017[50] NET017[51] NET017[52] NET017[53] NET017[54] 
+ NET017[55] NET017[56] NET017[57] NET017[58] NET017[59] NET017[60] NET017[61] 
+ NET017[62] NET017[63] NET017[64] NET017[65] NET017[66] NET017[67] NET017[68] 
+ NET017[69] NET017[70] NET017[71] NET017[72] NET017[73] NET017[74] NET017[75] 
+ NET017[76] NET017[77] NET017[78] NET017[79] NET017[80] NET017[81] NET017[82] 
+ NET017[83] NET017[84] NET017[85] NET017[86] NET017[87] NET017[88] NET017[89] 
+ NET017[90] NET017[91] NET017[92] NET017[93] NET017[94] NET017[95] NET017[96] 
+ NET017[97] NET017[98] NET017[99] NET017[100] NET017[101] NET017[102] 
+ NET017[103] NET017[104] NET017[105] NET017[106] NET017[107] NET017[108] 
+ NET017[109] NET017[110] NET017[111] NET017[112] NET017[113] NET017[114] 
+ NET017[115] NET017[116] NET017[117] NET017[118] NET017[119] NET017[120] 
+ NET017[121] NET017[122] NET017[123] NET017[124] NET017[125] NET017[126] 
+ NET017[127] NET017[128] NET017[129] NET017[130] NET017[131] NET017[132] 
+ NET017[133] NET017[134] NET017[135] NET017[136] NET017[137] NET017[138] 
+ NET017[139] NET017[140] NET017[141] NET017[142] NET017[143] NET017[144] 
+ NET017[145] NET017[146] NET017[147] NET017[148] NET017[149] NET017[150] 
+ NET017[151] NET017[152] NET017[153] NET017[154] NET017[155] NET017[156] 
+ NET017[157] NET017[158] NET017[159] NET017[160] NET017[161] NET017[162] 
+ NET017[163] NET017[164] NET017[165] NET017[166] NET017[167] NET017[168] 
+ NET017[169] NET017[170] NET017[171] NET017[172] NET017[173] NET017[174] 
+ NET017[175] NET017[176] NET017[177] NET017[178] NET017[179] NET017[180] 
+ NET017[181] NET017[182] NET017[183] NET017[184] NET017[185] NET017[186] 
+ NET017[187] NET017[188] NET017[189] NET017[190] NET017[191] NET017[192] 
+ NET017[193] NET017[194] NET017[195] NET017[196] NET017[197] NET017[198] 
+ NET017[199] NET017[200] NET017[201] NET017[202] NET017[203] NET017[204] 
+ NET017[205] NET017[206] NET017[207] NET017[208] NET017[209] NET017[210] 
+ NET017[211] NET017[212] NET017[213] NET017[214] NET017[215] NET017[216] 
+ NET017[217] NET017[218] NET017[219] NET017[220] NET017[221] NET017[222] 
+ NET017[223] NET017[224] NET017[225] NET017[226] NET017[227] NET017[228] 
+ NET017[229] NET017[230] NET017[231] NET017[232] NET017[233] NET017[234] 
+ NET017[235] NET017[236] NET017[237] NET017[238] NET017[239] NET017[240] 
+ NET017[241] NET017[242] NET017[243] NET017[244] NET017[245] NET017[246] 
+ NET017[247] NET017[248] NET017[249] NET017[250] NET017[251] 
+ S1AHSF400W40_MCB_252X4_SB_CHAR
XI36 NET8[0] NET8[1] NET8[2] NET8[3] NET7[0] NET7[1] NET7[2] NET7[3] NET9 
+ NET10 NET012[0] NET012[1] NET012[2] NET012[3] NET012[4] NET012[5] NET012[6] 
+ NET012[7] NET012[8] NET012[9] NET012[10] NET012[11] NET012[12] NET012[13] 
+ NET012[14] NET012[15] NET012[16] NET012[17] NET012[18] NET012[19] NET012[20] 
+ NET012[21] NET012[22] NET012[23] NET012[24] NET012[25] NET012[26] NET012[27] 
+ NET012[28] NET012[29] NET012[30] NET012[31] NET012[32] NET012[33] NET012[34] 
+ NET012[35] NET012[36] NET012[37] NET012[38] NET012[39] NET012[40] NET012[41] 
+ NET012[42] NET012[43] NET012[44] NET012[45] NET012[46] NET012[47] NET012[48] 
+ NET012[49] NET012[50] NET012[51] NET012[52] NET012[53] NET012[54] NET012[55] 
+ NET012[56] NET012[57] NET012[58] NET012[59] NET012[60] NET012[61] NET012[62] 
+ NET012[63] NET012[64] NET012[65] NET012[66] NET012[67] NET012[68] NET012[69] 
+ NET012[70] NET012[71] NET012[72] NET012[73] NET012[74] NET012[75] NET012[76] 
+ NET012[77] NET012[78] NET012[79] NET012[80] NET012[81] NET012[82] NET012[83] 
+ NET012[84] NET012[85] NET012[86] NET012[87] NET012[88] NET012[89] NET012[90] 
+ NET012[91] NET012[92] NET012[93] NET012[94] NET012[95] NET012[96] NET012[97] 
+ NET012[98] NET012[99] NET012[100] NET012[101] NET012[102] NET012[103] 
+ NET012[104] NET012[105] NET012[106] NET012[107] NET012[108] NET012[109] 
+ NET012[110] NET012[111] NET012[112] NET012[113] NET012[114] NET012[115] 
+ NET012[116] NET012[117] NET012[118] NET012[119] NET012[120] NET012[121] 
+ NET012[122] NET012[123] S1AHSF400W40_MCB_124X4_SB_CHAR
XI37 NET014[0] NET014[1] NET014[2] NET014[3] NET013[0] NET013[1] NET013[2] 
+ NET013[3] NET015 NET016 NET07[0] NET07[1] NET07[2] NET07[3] NET07[4] 
+ NET07[5] NET07[6] NET07[7] NET07[8] NET07[9] NET07[10] NET07[11] 
+ S1AHSF400W40_MCB_12X4_SB_CHAR
.ENDS

************************************************************************
* LIBRARY NAME: N65_LOGIC
* CELL NAME:    NAND3_BULK
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_NAND3_BULK A B C G GB P PB Y
*.PININFO A:I B:I C:I G:I GB:I P:I PB:I Y:O
M1 Y C P PB PCH L=LP3 W=WP3 M=1*FP3
M4 Y B P PB PCH L=LP2 W=WP2 M=1*FP2
M6 Y A P PB PCH L=LP1 W=WP1 M=1*FP1
M8 NET14 A G GB NCH L=LN1 W=WN1 M=1*FN1
M10 NET17 B NET14 GB NCH L=LN2 W=WN2 M=1*FN2
M12 Y C NET17 GB NCH L=LN3 W=WN3 M=1*FN3
.ENDS

************************************************************************
* LIBRARY NAME: N65_LOGIC
* CELL NAME:    AINV
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_AINV A G V Y
*.PININFO A:I G:I V:I Y:O
M1 Y A V V PCH L=LP W=WP M=1*FP
M3 Y A G G NCH L=LN W=WN M=1*FN
.ENDS

************************************************************************
* LIBRARY NAME: N65_LOGIC
* CELL NAME:    ANAND
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ANAND A B G V Y
*.PININFO A:I B:I G:I V:I Y:O
M1 Y B V V PCH L=LP2 W=WP2 M=1*FP2
M4 Y A V V PCH L=LP1 W=WP1 M=1*FP1
M6 NET9 A G G NCH L=LN1 W=WN1 M=1*FN1
M8 Y B NET9 G NCH L=LN2 W=WN2 M=1*FN2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    DOUT_M16_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_DOUT_M16_SB AWT AWTD BLEQ DL[0] DL[1] DLB[0] DLB[1] PD Q SAE2IO VDDHD 
+ VDDI VSSI YL[0] YL[1]
*.PININFO AWT:I AWTD:I BLEQ:I PD:I SAE2IO:I YL[0]:I YL[1]:I Q:O DL[0]:B 
*.PININFO DL[1]:B DLB[0]:B DLB[1]:B VDDHD:B VDDI:B VSSI:B
XI175 PREB SAE_OFF YL[0] VSSI VSSI VDDHD VDDHD PGB[0] S1AHSF400W40_NAND3_BULK FN3=1 
+ WN3=0.6U LN3=0.06U FN2=1 WN2=0.6U LN2=0.06U FN1=1 WN1=0.6U LN1=0.06U FP1=1 
+ WP1=0.3U LP1=0.06U FP2=1 WP2=0.3U LP2=0.06U FP3=1 WP3=0.3U LP3=0.06U M=1
XI176 PREB SAE_OFF YL[1] VSSI VSSI VDDHD VDDHD PGB[1] S1AHSF400W40_NAND3_BULK FN3=1 
+ WN3=0.6U LN3=0.06U FN2=1 WN2=0.6U LN2=0.06U FN1=1 WN1=0.6U LN1=0.06U FP1=1 
+ WP1=0.3U LP1=0.06U FP2=1 WP2=0.3U LP2=0.06U FP3=1 WP3=0.3U LP3=0.06U M=1
MM27 DLB_IN PGB[1] DLB[1] VDDI PCH L=60N W=1.2U M=1
MM2 VDDI PREB DL_IN VDDI PCH L=100N W=500N M=1
MM13 DL[1] PGB[1] DL_IN VDDI PCH L=60N W=1.2U M=1
MM31 DL[0] PGB[0] DL_IN VDDI PCH L=60N W=1.2U M=1
MM28 DLB_IN PGB[0] DLB[0] VDDI PCH L=60N W=1.2U M=1
MM1 DLB_IN PREB VDDI VDDI PCH L=100N W=500N M=1
MM20 NET0183 NET0249 VDDHD VDDHD PCH L=60N W=400N M=1
MM30 VDDHD DLB_IN NET0239 VDDHD PCH L=60N W=2U M=1
MM3 VDDI DLB_IN DL_IN VDDI PCH L=120.0N W=500N M=1
MP8 DL_IN PREB DLB_IN VDDI PCH L=120.0N W=500N M=2
MM17 NET0183 SAEBB QBB VDDHD PCH L=60N W=400N M=1
MM25 NET0187 SAEB QBB VDDHD PCH L=60N W=2U M=1
MP3 DLB_IN DL_IN VDDI VDDI PCH L=120.0N W=500N M=1
MM14 VDDHD DL_IN NET0187 VDDHD PCH L=60N W=2U M=1
MP10 VDDHD QBB Q VDDHD PCH L=60N W=750.0N M=2
MM10 PREB PD VSSI VSSI NCH L=60N W=600N M=1
MM11 SAE PD VSSI VSSI NCH L=60N W=600N M=1
MN2 NS SAE VSSI VSSI NCH L=80N W=750.0N M=4
MN0 NS DLB_IN DL_IN VSSI NCH L=180.0N W=750.0N M=4
MM4 DLB_IN DL_IN NS VSSI NCH L=180.0N W=750.0N M=4
MN5 Q QBB VSSI VSSI NCH L=60N W=800N M=1
MM5 Q PD VSSI VSSI NCH L=60N W=500N M=1
MM16 QBB SAEBB NET0263 VSSI NCH L=60N W=600N M=1
MM21 VSSI NET0249 NET0250 VSSI NCH L=60N W=400N M=1
MM18 QBB SAEB NET0250 VSSI NCH L=60N W=400N M=1
MM29 NET0239 DLB_IN VSSI VSSI NCH L=60N W=750.0N M=1
MM15 NET0263 DL_IN VSSI VSSI NCH L=60N W=750.0N M=1
XI161 SAEC VSSI VDDHD SAE S1AHSF400W40_AINV FN=1 WN=0.6U LN=0.06U FP=1 WP=0.8U LP=0.06U 
+ M=1
XI171 QBB VSSI VDDHD NET0249 S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 WP=0.2U 
+ LP=0.06U M=1
XI168 SAE VSSI VDDHD SAEB S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.6U LP=0.06U 
+ M=1
XI159 BLEQ VSSI VDDHD PREB S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.6U LP=0.06U 
+ M=1
XI170 SAEB VSSI VDDHD SAEBB S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.6U LP=0.06U 
+ M=1
XINV3 SAE_OFFB VSSI VDDHD SAE_OFF S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.3U 
+ LP=0.06U M=1
XI154 SAE_OFF SAE2IO VSSI VDDHD SAEC S1AHSF400W40_ANAND FN2=1 WN2=0.4U LN2=60N FN1=1 
+ WN1=0.4U LN1=60N FP1=1 WP1=0.3U LP1=60N FP2=1 WP2=0.3U LP2=60N M=1
XNAND2 DL_IN DLB_IN VSSI VDDHD SAE_OFFB S1AHSF400W40_ANAND FN2=1 WN2=0.2U LN2=0.06U FN1=1 
+ WN1=0.2U LN1=0.06U FP1=1 WP1=0.2U LP1=0.06U FP2=1 WP2=0.2U LP2=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65_LOGIC
* CELL NAME:    INV_BULK
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_INV_BULK A G GB P PB Y
*.PININFO A:I G:I GB:I P:I PB:I Y:O
M1 Y A P PB PCH L=LP W=WP M=1*FP
M3 Y A G GB NCH L=LN W=WN M=1*FN
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    DIN_M16_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_DIN_M16_SB AWTD BIST BWEB BWEBM CKD D DM VDDHD VSSI WC[0] WC[1] WT[0] 
+ WT[1] YL[0] YL[1]
*.PININFO BIST:I BWEB:I BWEBM:I CKD:I D:I DM:I YL[0]:I YL[1]:I AWTD:O WC[0]:O 
*.PININFO WC[1]:O WT[0]:O WT[1]:O VDDHD:B VSSI:B
XI353 CKD1B VSSI VSSI VDDHD VDDHD CKD2 S1AHSF400W40_INV_BULK FN=1 WN=0.6U LN=0.06U FP=1 
+ WP=1.2U LP=0.06U M=1
XI354 CKD VSSI VSSI VDDHD VDDHD CKD1B S1AHSF400W40_INV_BULK FN=1 WN=0.4U LN=0.06U FP=1 
+ WP=0.8U LP=0.06U M=1
XI76 GWB YL[0] VSSI VDDHD NET249 S1AHSF400W40_ANAND FN2=1 WN2=0.5U LN2=0.06U FN1=1 
+ WN1=0.5U LN1=0.06U FP1=1 WP1=0.5U LP1=0.06U FP2=1 WP2=0.5U LP2=0.06U M=1
XI281 GW YL[1] VSSI VDDHD NET239 S1AHSF400W40_ANAND FN2=1 WN2=0.5U LN2=0.06U FN1=1 
+ WN1=0.5U LN1=0.06U FP1=1 WP1=0.5U LP1=0.06U FP2=1 WP2=0.5U LP2=0.06U M=1
XI280 GWB YL[1] VSSI VDDHD NET234 S1AHSF400W40_ANAND FN2=1 WN2=0.5U LN2=0.06U FN1=1 
+ WN1=0.5U LN1=0.06U FP1=1 WP1=0.5U LP1=0.06U FP2=1 WP2=0.5U LP2=0.06U M=1
XI279 GW YL[0] VSSI VDDHD NET244 S1AHSF400W40_ANAND FN2=1 WN2=0.5U LN2=0.06U FN1=1 
+ WN1=0.5U LN1=0.06U FP1=1 WP1=0.5U LP1=0.06U FP2=1 WP2=0.5U LP2=0.06U M=1
MM70 BXL CKD1B Z16 VDDHD PCH L=120.0N W=600N M=1
MM72 DXL DXB Z9 VDDHD PCH L=120.0N W=600N M=1
MM73 DXL CKD1B Z6 VDDHD PCH L=120.0N W=600N M=1
MM76 BXL BXB Z13 VDDHD PCH L=120.0N W=600N M=1
MM66 DXL3B_AND BXL1B VDDHD VDDHD PCH L=60N W=500N M=2
MM61 DXL3B_AND DXL2 VDDHD VDDHD PCH L=60N W=500N M=2
MM62 VDDHD DXL1B Z6 VDDHD PCH L=120.0N W=600N M=1
MP10 DXL2_AND CKD2 VDDHD VDDHD PCH L=60N W=500N M=2
MP1 DXL3B_AND CKD2 VDDHD VDDHD PCH L=60N W=500N M=2
MM64 DXL2_AND DXL1B VDDHD VDDHD PCH L=60N W=500N M=2
MM65 DXL2_AND BXL1B VDDHD VDDHD PCH L=60N W=500N M=2
MM67 VDDHD CKD2 Z9 VDDHD PCH L=120.0N W=600N M=1
MM68 VDDHD CKD2 Z13 VDDHD PCH L=120.0N W=600N M=1
MM69 VDDHD BXL1B Z16 VDDHD PCH L=120.0N W=600N M=1
MM55 DXL DXB Z11 VSSI NCH L=120.0N W=300N M=1
MM54 VSSI CKD1B Z11 VSSI NCH L=120.0N W=300N M=1
MN33 DXL3B_AND DXL2 Z2 VSSI NCH L=60N W=1U M=2
MM50 BXL CKD2 Z14 VSSI NCH L=120.0N W=300N M=1
MN7 Z1 BXL1B VSSI VSSI NCH L=60N W=1U M=2
MN2 Z2 CKD2 Z1 VSSI NCH L=60N W=1U M=2
MM58 VSSI DXL1B Z7 VSSI NCH L=120.0N W=300N M=1
MM59 VSSI CKD1B Z15 VSSI NCH L=120.0N W=300N M=1
MM60 BXL BXB Z15 VSSI NCH L=120.0N W=300N M=1
MN1 DXL2_AND DXL1B Z2 VSSI NCH L=60N W=1U M=2
MM51 DXL CKD2 Z7 VSSI NCH L=120.0N W=300N M=1
MM49 VSSI BXL1B Z14 VSSI NCH L=120.0N W=300N M=1
XI358 NET0499 VSSI VDDHD WT[0] S1AHSF400W40_AINV FN=6 WN=0.8U LN=0.06U FP=6 WP=0.3U 
+ LP=0.06U M=1
XI360 NET0491 VSSI VDDHD WT[1] S1AHSF400W40_AINV FN=6 WN=0.8U LN=0.06U FP=6 WP=0.3U 
+ LP=0.06U M=1
XI359 NET0511 VSSI VDDHD WC[0] S1AHSF400W40_AINV FN=6 WN=0.8U LN=0.06U FP=6 WP=0.3U 
+ LP=0.06U M=1
XI276 NET244 VSSI VDDHD NET0511 S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U 
+ LP=0.06U M=1
XI277 NET234 VSSI VDDHD NET0491 S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U 
+ LP=0.06U M=1
XI347 DXL2_AND VSSI VDDHD GWB S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U LP=0.06U 
+ M=1
XI361 NET0487 VSSI VDDHD WC[1] S1AHSF400W40_AINV FN=6 WN=0.8U LN=0.06U FP=6 WP=0.3U 
+ LP=0.06U M=1
XI349 BXL VSSI VDDHD BXL1B S1AHSF400W40_AINV FN=2 WN=0.3U LN=0.06U FP=2 WP=0.6U LP=0.06U 
+ M=1
XI351 DXL VSSI VDDHD DXL1B S1AHSF400W40_AINV FN=2 WN=0.3U LN=0.06U FP=2 WP=0.6U LP=0.06U 
+ M=1
XINV01 D VSSI VDDHD DXB S1AHSF400W40_AINV FN=1 WN=0.3U LN=120N FP=1 WP=0.3U LP=120N M=1
XI254 DXL3B_AND VSSI VDDHD GW S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U LP=0.06U 
+ M=1
XI352 BWEB VSSI VDDHD BXB S1AHSF400W40_AINV FN=1 WN=0.3U LN=120N FP=1 WP=0.3U LP=120N M=1
XINV05 DXL1B VSSI VDDHD DXL2 S1AHSF400W40_AINV FN=2 WN=0.3U LN=0.06U FP=2 WP=0.6U 
+ LP=0.06U M=1
XINV1 NET249 VSSI VDDHD NET0499 S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U 
+ LP=0.06U M=1
XI278 NET239 VSSI VDDHD NET0487 S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U 
+ LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    PRECHARGE_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_PRECHARGE_SB BL BLB BLEQB VDDI
*.PININFO BLEQB:I BL:B BLB:B VDDI:B
MP17<0> BLB BLEQB VDDI VDDI PCH L=60N W=800N M=1
MP17<1> BLB BLEQB VDDI VDDI PCH L=60N W=800N M=1
MP17<2> BLB BLEQB VDDI VDDI PCH L=60N W=800N M=1
*MP5 BL BLEQB BLB VDDI PCH L=60N W=800N M=1
MP0<0> VDDI BLEQB BL VDDI PCH L=60N W=800N M=1
MP0<1> VDDI BLEQB BL VDDI PCH L=60N W=800N M=1
MP0<2> VDDI BLEQB BL VDDI PCH L=60N W=800N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    YPASS_M8_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_YPASS_M8_SB BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BLB[0] 
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLEQ DL DLB READ VDDI VSSI 
+ WC WRITE WT Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7]
*.PININFO BLEQ:I READ:I WRITE:I Y[0]:I Y[1]:I Y[2]:I Y[3]:I Y[4]:I Y[5]:I 
*.PININFO Y[6]:I Y[7]:I BL[0]:B BL[1]:B BL[2]:B BL[3]:B BL[4]:B BL[5]:B 
*.PININFO BL[6]:B BL[7]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B BLB[4]:B 
*.PININFO BLB[5]:B BLB[6]:B BLB[7]:B DL:B DLB:B VDDI:B VSSI:B WC:B WT:B
MN1<0> NET88[0] WRITE VSSI VSSI NCH L=60N W=200N M=1
MN1<1> NET88[1] WRITE VSSI VSSI NCH L=60N W=200N M=1
MN1<2> NET88[2] WRITE VSSI VSSI NCH L=60N W=200N M=1
MN1<3> NET88[3] WRITE VSSI VSSI NCH L=60N W=200N M=1
MN1<4> NET88[4] WRITE VSSI VSSI NCH L=60N W=200N M=1
MN1<5> NET88[5] WRITE VSSI VSSI NCH L=60N W=200N M=1
MN1<6> NET88[6] WRITE VSSI VSSI NCH L=60N W=200N M=1
MN1<7> NET88[7] WRITE VSSI VSSI NCH L=60N W=200N M=1
MN31<0> BL[0] Y_WRITE[0] WT VSSI NCH L=60N W=1.6U M=1
MN31<1> BL[1] Y_WRITE[1] WT VSSI NCH L=60N W=1.6U M=1
MN31<2> BL[2] Y_WRITE[2] WT VSSI NCH L=60N W=1.6U M=1
MN31<3> BL[3] Y_WRITE[3] WT VSSI NCH L=60N W=1.6U M=1
MN31<4> BL[4] Y_WRITE[4] WT VSSI NCH L=60N W=1.6U M=1
MN31<5> BL[5] Y_WRITE[5] WT VSSI NCH L=60N W=1.6U M=1
MN31<6> BL[6] Y_WRITE[6] WT VSSI NCH L=60N W=1.6U M=1
MN31<7> BL[7] Y_WRITE[7] WT VSSI NCH L=60N W=1.6U M=1
MN13<0> NET84[0] READ VSSI VSSI NCH L=60N W=200N M=1
MN13<1> NET84[1] READ VSSI VSSI NCH L=60N W=200N M=1
MN13<2> NET84[2] READ VSSI VSSI NCH L=60N W=200N M=1
MN13<3> NET84[3] READ VSSI VSSI NCH L=60N W=200N M=1
MN13<4> NET84[4] READ VSSI VSSI NCH L=60N W=200N M=1
MN13<5> NET84[5] READ VSSI VSSI NCH L=60N W=200N M=1
MN13<6> NET84[6] READ VSSI VSSI NCH L=60N W=200N M=1
MN13<7> NET84[7] READ VSSI VSSI NCH L=60N W=200N M=1
MN18<0> BLB[0] Y_WRITE[0] WC VSSI NCH L=60N W=1.6U M=1
MN18<1> BLB[1] Y_WRITE[1] WC VSSI NCH L=60N W=1.6U M=1
MN18<2> BLB[2] Y_WRITE[2] WC VSSI NCH L=60N W=1.6U M=1
MN18<3> BLB[3] Y_WRITE[3] WC VSSI NCH L=60N W=1.6U M=1
MN18<4> BLB[4] Y_WRITE[4] WC VSSI NCH L=60N W=1.6U M=1
MN18<5> BLB[5] Y_WRITE[5] WC VSSI NCH L=60N W=1.6U M=1
MN18<6> BLB[6] Y_WRITE[6] WC VSSI NCH L=60N W=1.6U M=1
MN18<7> BLB[7] Y_WRITE[7] WC VSSI NCH L=60N W=1.6U M=1
MP29<0> YB_WRITE[0] WRITE VDDI VDDI PCH L=60N W=200N M=1
MP29<1> YB_WRITE[1] WRITE VDDI VDDI PCH L=60N W=200N M=1
MP29<2> YB_WRITE[2] WRITE VDDI VDDI PCH L=60N W=200N M=1
MP29<3> YB_WRITE[3] WRITE VDDI VDDI PCH L=60N W=200N M=1
MP29<4> YB_WRITE[4] WRITE VDDI VDDI PCH L=60N W=200N M=1
MP29<5> YB_WRITE[5] WRITE VDDI VDDI PCH L=60N W=200N M=1
MP29<6> YB_WRITE[6] WRITE VDDI VDDI PCH L=60N W=200N M=1
MP29<7> YB_WRITE[7] WRITE VDDI VDDI PCH L=60N W=200N M=1
MP22 VDDI BLEQB DL VDDI PCH L=60N W=200N M=1
MP0<0> DL YB_READ[0] BL[0] VDDI PCH L=60N W=800N M=1
MP0<1> DL YB_READ[1] BL[1] VDDI PCH L=60N W=800N M=1
MP0<2> DL YB_READ[2] BL[2] VDDI PCH L=60N W=800N M=1
MP0<3> DL YB_READ[3] BL[3] VDDI PCH L=60N W=800N M=1
MP0<4> DL YB_READ[4] BL[4] VDDI PCH L=60N W=800N M=1
MP0<5> DL YB_READ[5] BL[5] VDDI PCH L=60N W=800N M=1
MP0<6> DL YB_READ[6] BL[6] VDDI PCH L=60N W=800N M=1
MP0<7> DL YB_READ[7] BL[7] VDDI PCH L=60N W=800N M=1
MP3 DLB BLEQB VDDI VDDI PCH L=60N W=200N M=1
MP17<0> YB_READ[0] READ VDDI VDDI PCH L=60N W=200N M=1
MP17<1> YB_READ[1] READ VDDI VDDI PCH L=60N W=200N M=1
MP17<2> YB_READ[2] READ VDDI VDDI PCH L=60N W=200N M=1
MP17<3> YB_READ[3] READ VDDI VDDI PCH L=60N W=200N M=1
MP17<4> YB_READ[4] READ VDDI VDDI PCH L=60N W=200N M=1
MP17<5> YB_READ[5] READ VDDI VDDI PCH L=60N W=200N M=1
MP17<6> YB_READ[6] READ VDDI VDDI PCH L=60N W=200N M=1
MP17<7> YB_READ[7] READ VDDI VDDI PCH L=60N W=200N M=1
MP10<0> DLB YB_READ[0] BLB[0] VDDI PCH L=60N W=800N M=1
MP10<1> DLB YB_READ[1] BLB[1] VDDI PCH L=60N W=800N M=1
MP10<2> DLB YB_READ[2] BLB[2] VDDI PCH L=60N W=800N M=1
MP10<3> DLB YB_READ[3] BLB[3] VDDI PCH L=60N W=800N M=1
MP10<4> DLB YB_READ[4] BLB[4] VDDI PCH L=60N W=800N M=1
MP10<5> DLB YB_READ[5] BLB[5] VDDI PCH L=60N W=800N M=1
MP10<6> DLB YB_READ[6] BLB[6] VDDI PCH L=60N W=800N M=1
MP10<7> DLB YB_READ[7] BLB[7] VDDI PCH L=60N W=800N M=1
XI252<0> Y[0] NET88[0] VSSI VDDI VDDI YB_WRITE[0] S1AHSF400W40_INV_BULK FN=1 WN=0.2U 
+ LN=0.06U FP=1 WP=0.2U LP=0.06U M=1
XI252<1> Y[1] NET88[1] VSSI VDDI VDDI YB_WRITE[1] S1AHSF400W40_INV_BULK FN=1 WN=0.2U 
+ LN=0.06U FP=1 WP=0.2U LP=0.06U M=1
XI252<2> Y[2] NET88[2] VSSI VDDI VDDI YB_WRITE[2] S1AHSF400W40_INV_BULK FN=1 WN=0.2U 
+ LN=0.06U FP=1 WP=0.2U LP=0.06U M=1
XI252<3> Y[3] NET88[3] VSSI VDDI VDDI YB_WRITE[3] S1AHSF400W40_INV_BULK FN=1 WN=0.2U 
+ LN=0.06U FP=1 WP=0.2U LP=0.06U M=1
XI252<4> Y[4] NET88[4] VSSI VDDI VDDI YB_WRITE[4] S1AHSF400W40_INV_BULK FN=1 WN=0.2U 
+ LN=0.06U FP=1 WP=0.2U LP=0.06U M=1
XI252<5> Y[5] NET88[5] VSSI VDDI VDDI YB_WRITE[5] S1AHSF400W40_INV_BULK FN=1 WN=0.2U 
+ LN=0.06U FP=1 WP=0.2U LP=0.06U M=1
XI252<6> Y[6] NET88[6] VSSI VDDI VDDI YB_WRITE[6] S1AHSF400W40_INV_BULK FN=1 WN=0.2U 
+ LN=0.06U FP=1 WP=0.2U LP=0.06U M=1
XI252<7> Y[7] NET88[7] VSSI VDDI VDDI YB_WRITE[7] S1AHSF400W40_INV_BULK FN=1 WN=0.2U 
+ LN=0.06U FP=1 WP=0.2U LP=0.06U M=1
XI249<0> Y[0] NET84[0] VSSI VDDI VDDI YB_READ[0] S1AHSF400W40_INV_BULK FN=1 WN=0.2U 
+ LN=0.06U FP=1 WP=0.2U LP=0.06U M=1
XI249<1> Y[1] NET84[1] VSSI VDDI VDDI YB_READ[1] S1AHSF400W40_INV_BULK FN=1 WN=0.2U 
+ LN=0.06U FP=1 WP=0.2U LP=0.06U M=1
XI249<2> Y[2] NET84[2] VSSI VDDI VDDI YB_READ[2] S1AHSF400W40_INV_BULK FN=1 WN=0.2U 
+ LN=0.06U FP=1 WP=0.2U LP=0.06U M=1
XI249<3> Y[3] NET84[3] VSSI VDDI VDDI YB_READ[3] S1AHSF400W40_INV_BULK FN=1 WN=0.2U 
+ LN=0.06U FP=1 WP=0.2U LP=0.06U M=1
XI249<4> Y[4] NET84[4] VSSI VDDI VDDI YB_READ[4] S1AHSF400W40_INV_BULK FN=1 WN=0.2U 
+ LN=0.06U FP=1 WP=0.2U LP=0.06U M=1
XI249<5> Y[5] NET84[5] VSSI VDDI VDDI YB_READ[5] S1AHSF400W40_INV_BULK FN=1 WN=0.2U 
+ LN=0.06U FP=1 WP=0.2U LP=0.06U M=1
XI249<6> Y[6] NET84[6] VSSI VDDI VDDI YB_READ[6] S1AHSF400W40_INV_BULK FN=1 WN=0.2U 
+ LN=0.06U FP=1 WP=0.2U LP=0.06U M=1
XI249<7> Y[7] NET84[7] VSSI VDDI VDDI YB_READ[7] S1AHSF400W40_INV_BULK FN=1 WN=0.2U 
+ LN=0.06U FP=1 WP=0.2U LP=0.06U M=1
XPRECHARGE<0> BLB[0] BL[0] BLEQB VDDI S1AHSF400W40_PRECHARGE_SB
XPRECHARGE<1> BLB[1] BL[1] BLEQB VDDI S1AHSF400W40_PRECHARGE_SB
XPRECHARGE<2> BLB[2] BL[2] BLEQB VDDI S1AHSF400W40_PRECHARGE_SB
XPRECHARGE<3> BLB[3] BL[3] BLEQB VDDI S1AHSF400W40_PRECHARGE_SB
XPRECHARGE<4> BLB[4] BL[4] BLEQB VDDI S1AHSF400W40_PRECHARGE_SB
XPRECHARGE<5> BLB[5] BL[5] BLEQB VDDI S1AHSF400W40_PRECHARGE_SB
XPRECHARGE<6> BLB[6] BL[6] BLEQB VDDI S1AHSF400W40_PRECHARGE_SB
XPRECHARGE<7> BLB[7] BL[7] BLEQB VDDI S1AHSF400W40_PRECHARGE_SB
XI214<0> YB_WRITE[0] VSSI VDDI Y_WRITE[0] S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 
+ WP=0.2U LP=0.06U M=1
XI214<1> YB_WRITE[1] VSSI VDDI Y_WRITE[1] S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 
+ WP=0.2U LP=0.06U M=1
XI214<2> YB_WRITE[2] VSSI VDDI Y_WRITE[2] S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 
+ WP=0.2U LP=0.06U M=1
XI214<3> YB_WRITE[3] VSSI VDDI Y_WRITE[3] S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 
+ WP=0.2U LP=0.06U M=1
XI214<4> YB_WRITE[4] VSSI VDDI Y_WRITE[4] S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 
+ WP=0.2U LP=0.06U M=1
XI214<5> YB_WRITE[5] VSSI VDDI Y_WRITE[5] S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 
+ WP=0.2U LP=0.06U M=1
XI214<6> YB_WRITE[6] VSSI VDDI Y_WRITE[6] S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 
+ WP=0.2U LP=0.06U M=1
XI214<7> YB_WRITE[7] VSSI VDDI Y_WRITE[7] S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 
+ WP=0.2U LP=0.06U M=1
XINV0 BLEQ VSSI VDDI BLEQB S1AHSF400W40_AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=1.6U LP=0.06U 
+ M=2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MIO_M16_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MIO_M16_SB AWT2 BIST2IO BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] 
+ BL[7] BL[8] BL[9] BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BLB[0] BLB[1] 
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] 
+ BLB[12] BLB[13] BLB[14] BLB[15] BLEQ BWEB BWEBM CKD D DM PD_BUF Q RE SAE 
+ VDDHD VDDI VSSI WE Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7] YL[0] YL[1]
*.PININFO AWT2:I BIST2IO:I BLEQ:I BWEB:I BWEBM:I CKD:I D:I DM:I PD_BUF:I RE:I 
*.PININFO SAE:I WE:I Y[0]:I Y[1]:I Y[2]:I Y[3]:I Y[4]:I Y[5]:I Y[6]:I Y[7]:I 
*.PININFO YL[0]:I YL[1]:I Q:O BL[0]:B BL[1]:B BL[2]:B BL[3]:B BL[4]:B BL[5]:B 
*.PININFO BL[6]:B BL[7]:B BL[8]:B BL[9]:B BL[10]:B BL[11]:B BL[12]:B BL[13]:B 
*.PININFO BL[14]:B BL[15]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B BLB[4]:B 
*.PININFO BLB[5]:B BLB[6]:B BLB[7]:B BLB[8]:B BLB[9]:B BLB[10]:B BLB[11]:B 
*.PININFO BLB[12]:B BLB[13]:B BLB[14]:B BLB[15]:B VDDHD:B VDDI:B VSSI:B
MP10 VDDHD PD_BUF VDDI VDDI PCH L=65.0N W=2.5U M=2
MM0 VDDHD PD_BUF VDDI VDDI PCH L=60N W=1U M=10
XDOUT AWT2 AWTD BLEQI DL[0] DL[1] DLB[0] DLB[1] PD_BUF Q SAE VDDHD VDDI VSSI 
+ YL[0] YL[1] S1AHSF400W40_DOUT_M16_SB
XDIN AWTD BIST2IO BWEB BWEBM CKD D DM VDDHD VSSI WC[0] WC[1] WT[0] WT[1] YL[0] 
+ YL[1] S1AHSF400W40_DIN_M16_SB
XYPASS BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BLB[0] BLB[1] BLB[2] 
+ BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLEQI DL[0] DLB[0] REI VDDI VSSI WC[0] 
+ WEI WT[0] Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7] S1AHSF400W40_YPASS_M8_SB
XYPASS_1 BL[8] BL[9] BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BLB[8] BLB[9] 
+ BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15] BLEQI DL[1] DLB[1] REI VDDI 
+ VSSI WC[1] WEI WT[1] Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7] S1AHSF400W40_YPASS_M8_SB
XI184 BLEQ VSSI VDDI BLEQI S1AHSF400W40_AINV FN=4 WN=0.2U LN=0.06U FP=4 WP=0.4U LP=0.06U 
+ M=1
XI213 WE VSSI VDDI NET280 S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 WP=0.4U LP=0.06U 
+ M=1
XI214 NET280 VSSI VDDI WEI S1AHSF400W40_AINV FN=1 WN=0.4U LN=0.06U FP=1 WP=0.8U LP=0.06U 
+ M=1
XI215 NET268 VSSI VDDI REI S1AHSF400W40_AINV FN=1 WN=0.4U LN=0.06U FP=1 WP=0.8U LP=0.06U 
+ M=1
XI216 RE VSSI VDDI NET268 S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 WP=0.4U LP=0.06U 
+ M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    DOUT_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_DOUT_SB AWT AWTD BLEQ DL DLB PD Q SAE2IO VDDHD VDDI VSSI
*.PININFO AWT:I AWTD:I BLEQ:I PD:I SAE2IO:I Q:O DL:B DLB:B VDDHD:B VDDI:B 
*.PININFO VSSI:B
XNAND2 DL_IN DLB_IN VSSI VDDHD SAE_OFFB S1AHSF400W40_ANAND FN2=1 WN2=0.2U LN2=0.06U FN1=1 
+ WN1=0.2U LN1=0.06U FP1=1 WP1=0.2U LP1=0.06U FP2=1 WP2=0.2U LP2=0.06U M=1
XI160 PREB SAE_OFF VSSI VDDHD PGB S1AHSF400W40_ANAND FN2=1 WN2=0.4U LN2=60N FN1=1 
+ WN1=0.4U LN1=60N FP1=1 WP1=0.3U LP1=60N FP2=1 WP2=0.3U LP2=60N M=1
XI154 SAE_OFF SAE2IO VSSI VDDHD SAEC S1AHSF400W40_ANAND FN2=1 WN2=0.4U LN2=60N FN1=1 
+ WN1=0.4U LN1=60N FP1=1 WP1=0.3U LP1=60N FP2=1 WP2=0.3U LP2=60N M=1
XI159 BLEQ VSSI VDDHD PREB S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.6U LP=0.06U 
+ M=1
XINV3 SAE_OFFB VSSI VDDHD SAE_OFF S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.3U 
+ LP=0.06U M=1
XI161 SAEC VSSI VDDHD SAE S1AHSF400W40_AINV FN=1 WN=0.6U LN=0.06U FP=1 WP=0.8U LP=0.06U 
+ M=1
XI163 QBB VSSI VDDHD NET243 S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 WP=0.2U LP=0.06U 
+ M=1
XI165 SAEB VSSI VDDHD SAEBB S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.6U LP=0.06U 
+ M=1
XI166 SAE VSSI VDDHD SAEB S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.6U LP=0.06U 
+ M=1
MM29 NET249 DLB_IN VSSI VSSI NCH L=60N W=750.0N M=1
MN5 Q QBB VSSI VSSI NCH L=60N W=800N M=1
MM10 PREB PD VSSI VSSI NCH L=60N W=600N M=1
MM18 QBB SAEB NET244 VSSI NCH L=60N W=400N M=1
MM21 VSSI NET243 NET244 VSSI NCH L=60N W=400N M=1
MM16 QBB SAEBB NET205 VSSI NCH L=60N W=600N M=1
MM15 NET205 DL_IN VSSI VSSI NCH L=60N W=750.0N M=1
MM11 SAE PD VSSI VSSI NCH L=60N W=600N M=1
MN0 NS DLB_IN DL_IN VSSI NCH L=180.0N W=750.0N M=4
MM4 DLB_IN DL_IN NS VSSI NCH L=180.0N W=750.0N M=4
MN2 NS SAE VSSI VSSI NCH L=80N W=750.0N M=4
MM5 Q PD VSSI VSSI NCH L=60N W=500N M=1
MM14 VDDHD DL_IN NET293 VDDHD PCH L=60N W=2U M=1
MM25 NET293 SAEB QBB VDDHD PCH L=60N W=2U M=1
MM20 NET297 NET243 VDDHD VDDHD PCH L=60N W=400N M=1
MM30 VDDHD DLB_IN NET249 VDDHD PCH L=60N W=2U M=1
MP7 DLB_IN PGB DLB VDDI PCH L=60N W=1.2U M=1
MP3 DLB_IN DL_IN VDDI VDDI PCH L=120.0N W=500N M=1
MM1 DLB_IN PREB VDDI VDDI PCH L=100N W=500N M=1
MP8 DL_IN PREB DLB_IN VDDI PCH L=120.0N W=500N M=2
MM3 VDDI DLB_IN DL_IN VDDI PCH L=120.0N W=500N M=1
MM0 DL PGB DL_IN VDDI PCH L=60N W=1.2U M=1
MM2 VDDI PREB DL_IN VDDI PCH L=100N W=500N M=1
MP10 VDDHD QBB Q VDDHD PCH L=60N W=750.0N M=2
MM17 NET297 SAEBB QBB VDDHD PCH L=60N W=400N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    DIN_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_DIN_SB AWTD BIST BWEB BWEBM CKD D DM VDDHD VSSI WC WT
*.PININFO BIST:I BWEB:I BWEBM:I CKD:I D:I DM:I AWTD:O WC:O WT:O VDDHD:B VSSI:B
XINV01 D VSSI VDDHD DXB S1AHSF400W40_AINV FN=1 WN=0.3U LN=120N FP=1 WP=0.3U LP=120N M=1
XI317 GWB VSSI VDDHD WT S1AHSF400W40_AINV FN=6 WN=0.8U LN=0.06U FP=6 WP=0.4U LP=0.06U M=1
XI319 BXL VSSI VDDHD BXL1B S1AHSF400W40_AINV FN=2 WN=0.3U LN=0.06U FP=2 WP=0.6U LP=0.06U 
+ M=1
XI318 DXL VSSI VDDHD DXL1B S1AHSF400W40_AINV FN=2 WN=0.3U LN=0.06U FP=2 WP=0.6U LP=0.06U 
+ M=1
XI254 DXL3B_AND VSSI VDDHD GW S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U LP=0.06U 
+ M=1
XI267 DXL2_AND VSSI VDDHD GWB S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U LP=0.06U 
+ M=1
XINV07 GW VSSI VDDHD WC S1AHSF400W40_AINV FN=6 WN=0.8U LN=0.06U FP=6 WP=0.4U LP=0.06U M=1
XINV05 DXL1B VSSI VDDHD DXL2 S1AHSF400W40_AINV FN=2 WN=0.3U LN=0.06U FP=2 WP=0.6U 
+ LP=0.06U M=1
XI352 BWEB VSSI VDDHD BXB S1AHSF400W40_AINV FN=1 WN=0.3U LN=120N FP=1 WP=0.3U LP=120N M=1
MM44 VSSI BXL1B Z14 VSSI NCH L=120.0N W=300N M=1
MM45 BXL CKD2 Z14 VSSI NCH L=120.0N W=300N M=1
MN7 Z1 BXL1B VSSI VSSI NCH L=60N W=1U M=2
MN1 DXL2_AND DXL1B Z2 VSSI NCH L=60N W=1U M=2
MM35 DXL CKD2 Z7 VSSI NCH L=120.0N W=300N M=1
MN33 DXL3B_AND DXL2 Z2 VSSI NCH L=60N W=1U M=2
MM36 VSSI CKD1B Z11 VSSI NCH L=120.0N W=300N M=1
MM34 DXL DXB Z11 VSSI NCH L=120.0N W=300N M=1
MN2 Z2 CKD2 Z1 VSSI NCH L=60N W=1U M=2
MM37 VSSI DXL1B Z7 VSSI NCH L=120.0N W=300N M=1
MM43 VSSI CKD1B Z15 VSSI NCH L=120.0N W=300N M=1
MM42 BXL BXB Z15 VSSI NCH L=120.0N W=300N M=1
MM51 DXL3B_AND DXL2 VDDHD VDDHD PCH L=60N W=500N M=2
MM28 VDDHD DXL1B Z6 VDDHD PCH L=120.0N W=600N M=1
MP10 DXL2_AND CKD2 VDDHD VDDHD PCH L=60N W=500N M=2
MP1 DXL3B_AND CKD2 VDDHD VDDHD PCH L=60N W=500N M=2
MM52 DXL2_AND DXL1B VDDHD VDDHD PCH L=60N W=500N M=2
MM53 DXL2_AND BXL1B VDDHD VDDHD PCH L=60N W=500N M=2
MM54 DXL3B_AND BXL1B VDDHD VDDHD PCH L=60N W=500N M=2
MM26 VDDHD CKD2 Z9 VDDHD PCH L=120.0N W=600N M=1
MM38 VDDHD CKD2 Z13 VDDHD PCH L=120.0N W=600N M=1
MM39 VDDHD BXL1B Z16 VDDHD PCH L=120.0N W=600N M=1
MM40 BXL CKD1B Z16 VDDHD PCH L=120.0N W=600N M=1
MM27 DXL DXB Z9 VDDHD PCH L=120.0N W=600N M=1
MM29 DXL CKD1B Z6 VDDHD PCH L=120.0N W=600N M=1
MM41 BXL BXB Z13 VDDHD PCH L=120.0N W=600N M=1
XI324 CKD1B VSSI VSSI VDDHD VDDHD CKD2 S1AHSF400W40_INV_BULK FN=1 WN=0.6U LN=0.06U FP=1 
+ WP=1.2U LP=0.06U M=1
XI323 CKD VSSI VSSI VDDHD VDDHD CKD1B S1AHSF400W40_INV_BULK FN=1 WN=0.4U LN=0.06U FP=1 
+ WP=0.8U LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MIO_M8_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MIO_M8_SB AWT2 BIST2IO BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] 
+ BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLEQ BWEB BWEBM CKD 
+ D DM PD_BUF Q RE SAE VDDHD VDDI VSSI WE Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] 
+ Y[7]
*.PININFO AWT2:I BIST2IO:I BLEQ:I BWEB:I BWEBM:I CKD:I D:I DM:I PD_BUF:I RE:I 
*.PININFO SAE:I WE:I Y[0]:I Y[1]:I Y[2]:I Y[3]:I Y[4]:I Y[5]:I Y[6]:I Y[7]:I 
*.PININFO Q:O BL[0]:B BL[1]:B BL[2]:B BL[3]:B BL[4]:B BL[5]:B BL[6]:B BL[7]:B 
*.PININFO BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B BLB[4]:B BLB[5]:B BLB[6]:B 
*.PININFO BLB[7]:B VDDHD:B VDDI:B VSSI:B
MP10 VDDHD PD_BUF VDDI VDDI PCH L=65.0N W=2.5U M=2
XDOUT AWT2 AWTD BLEQI DL DLB PD_BUF Q SAE VDDHD VDDI VSSI S1AHSF400W40_DOUT_SB
XDIN AWTD BIST2IO BWEB BWEBM CKD D DM VDDHD VSSI WC WT S1AHSF400W40_DIN_SB
XYPASS BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BLB[0] BLB[1] BLB[2] 
+ BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLEQI DL DLB REI VDDI VSSI WC WEI WT Y[0] 
+ Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7] S1AHSF400W40_YPASS_M8_SB
XI216 RE VSSI VDDI NET101 S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 WP=0.4U LP=0.06U 
+ M=1
XI215 NET101 VSSI VDDI REI S1AHSF400W40_AINV FN=1 WN=0.4U LN=0.06U FP=1 WP=0.8U LP=0.06U 
+ M=1
XI213 WE VSSI VDDI NET89 S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 WP=0.4U LP=0.06U M=1
XI184 BLEQ VSSI VDDI BLEQI S1AHSF400W40_AINV FN=2 WN=0.25U LN=0.06U FP=2 WP=0.5U LP=0.06U 
+ M=1
XI214 NET89 VSSI VDDI WEI S1AHSF400W40_AINV FN=1 WN=0.4U LN=0.06U FP=1 WP=0.8U LP=0.06U 
+ M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    YPASS_M4_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_YPASS_M4_SB BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] BLEQ 
+ DL DLB READ VDDI VSSI WC WRITE WT Y[0] Y[1] Y[2] Y[3]
*.PININFO BLEQ:I READ:I WRITE:I Y[0]:I Y[1]:I Y[2]:I Y[3]:I BL[0]:B BL[1]:B 
*.PININFO BL[2]:B BL[3]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B DL:B DLB:B 
*.PININFO VDDI:B VSSI:B WC:B WT:B
XPRECHARGE<0> BL[0] BLB[0] BLEQB VDDI S1AHSF400W40_PRECHARGE_SB
XPRECHARGE<1> BL[1] BLB[1] BLEQB VDDI S1AHSF400W40_PRECHARGE_SB
XPRECHARGE<2> BL[2] BLB[2] BLEQB VDDI S1AHSF400W40_PRECHARGE_SB
XPRECHARGE<3> BL[3] BLB[3] BLEQB VDDI S1AHSF400W40_PRECHARGE_SB
XINV0 BLEQ VSSI VDDI BLEQB S1AHSF400W40_AINV FN=1 WN=0.75U LN=0.06U FP=1 WP=1.55U 
+ LP=0.06U M=1
XI238<0> YB_WRITE[0] VSSI VDDI Y_WRITE[0] S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 
+ WP=0.2U LP=0.06U M=1
XI238<1> YB_WRITE[1] VSSI VDDI Y_WRITE[1] S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 
+ WP=0.2U LP=0.06U M=1
XI238<2> YB_WRITE[2] VSSI VDDI Y_WRITE[2] S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 
+ WP=0.2U LP=0.06U M=1
XI238<3> YB_WRITE[3] VSSI VDDI Y_WRITE[3] S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 
+ WP=0.2U LP=0.06U M=1
MN31<0> BL[0] Y_WRITE[0] WT VSSI NCH L=60N W=1.6U M=1
MN31<1> BL[1] Y_WRITE[1] WT VSSI NCH L=60N W=1.6U M=1
MN31<2> BL[2] Y_WRITE[2] WT VSSI NCH L=60N W=1.6U M=1
MN31<3> BL[3] Y_WRITE[3] WT VSSI NCH L=60N W=1.6U M=1
MN30<0> BLB[0] Y_WRITE[0] WC VSSI NCH L=60N W=1.6U M=1
MN30<1> BLB[1] Y_WRITE[1] WC VSSI NCH L=60N W=1.6U M=1
MN30<2> BLB[2] Y_WRITE[2] WC VSSI NCH L=60N W=1.6U M=1
MN30<3> BLB[3] Y_WRITE[3] WC VSSI NCH L=60N W=1.6U M=1
MN13<0> NET177[0] READ VSSI VSSI NCH L=60N W=200N M=1
MN13<1> NET177[1] READ VSSI VSSI NCH L=60N W=200N M=1
MN13<2> NET177[2] READ VSSI VSSI NCH L=60N W=200N M=1
MN13<3> NET177[3] READ VSSI VSSI NCH L=60N W=200N M=1
MM1<0> NET173[0] WRITE VSSI VSSI NCH L=60N W=200N M=1
MM1<1> NET173[1] WRITE VSSI VSSI NCH L=60N W=200N M=1
MM1<2> NET173[2] WRITE VSSI VSSI NCH L=60N W=200N M=1
MM1<3> NET173[3] WRITE VSSI VSSI NCH L=60N W=200N M=1
MP0 VDDI BLEQB DL VDDI PCH L=60N W=200N M=1
MP1<0> DL YB[0] BL[0] VDDI PCH L=60N W=800N M=1
MP1<1> DL YB[1] BL[1] VDDI PCH L=60N W=800N M=1
MP1<2> DL YB[2] BL[2] VDDI PCH L=60N W=800N M=1
MP1<3> DL YB[3] BL[3] VDDI PCH L=60N W=800N M=1
MP17<0> YB[0] READ VDDI VDDI PCH L=60N W=200N M=1
MP17<1> YB[1] READ VDDI VDDI PCH L=60N W=200N M=1
MP17<2> YB[2] READ VDDI VDDI PCH L=60N W=200N M=1
MP17<3> YB[3] READ VDDI VDDI PCH L=60N W=200N M=1
MM0<0> YB_WRITE[0] WRITE VDDI VDDI PCH L=60N W=200N M=1
MM0<1> YB_WRITE[1] WRITE VDDI VDDI PCH L=60N W=200N M=1
MM0<2> YB_WRITE[2] WRITE VDDI VDDI PCH L=60N W=200N M=1
MM0<3> YB_WRITE[3] WRITE VDDI VDDI PCH L=60N W=200N M=1
MP10<0> DLB YB[0] BLB[0] VDDI PCH L=60N W=800N M=1
MP10<1> DLB YB[1] BLB[1] VDDI PCH L=60N W=800N M=1
MP10<2> DLB YB[2] BLB[2] VDDI PCH L=60N W=800N M=1
MP10<3> DLB YB[3] BLB[3] VDDI PCH L=60N W=800N M=1
MP2 DLB BLEQB VDDI VDDI PCH L=60N W=200N M=1
XI281<0> Y[0] NET173[0] VSSI VDDI VDDI YB_WRITE[0] S1AHSF400W40_INV_BULK FN=1 WN=0.2U 
+ LN=0.06U FP=1 WP=0.2U LP=0.06U M=1
XI281<1> Y[1] NET173[1] VSSI VDDI VDDI YB_WRITE[1] S1AHSF400W40_INV_BULK FN=1 WN=0.2U 
+ LN=0.06U FP=1 WP=0.2U LP=0.06U M=1
XI281<2> Y[2] NET173[2] VSSI VDDI VDDI YB_WRITE[2] S1AHSF400W40_INV_BULK FN=1 WN=0.2U 
+ LN=0.06U FP=1 WP=0.2U LP=0.06U M=1
XI281<3> Y[3] NET173[3] VSSI VDDI VDDI YB_WRITE[3] S1AHSF400W40_INV_BULK FN=1 WN=0.2U 
+ LN=0.06U FP=1 WP=0.2U LP=0.06U M=1
XI249<0> Y[0] NET177[0] VSSI VDDI VDDI YB[0] S1AHSF400W40_INV_BULK FN=1 WN=0.2U LN=0.06U 
+ FP=1 WP=0.2U LP=0.06U M=1
XI249<1> Y[1] NET177[1] VSSI VDDI VDDI YB[1] S1AHSF400W40_INV_BULK FN=1 WN=0.2U LN=0.06U 
+ FP=1 WP=0.2U LP=0.06U M=1
XI249<2> Y[2] NET177[2] VSSI VDDI VDDI YB[2] S1AHSF400W40_INV_BULK FN=1 WN=0.2U LN=0.06U 
+ FP=1 WP=0.2U LP=0.06U M=1
XI249<3> Y[3] NET177[3] VSSI VDDI VDDI YB[3] S1AHSF400W40_INV_BULK FN=1 WN=0.2U LN=0.06U 
+ FP=1 WP=0.2U LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MIO_M4_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MIO_M4_SB AWT2 BIST2IO BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] 
+ BLB[3] BLEQ BWEB BWEBM CKD D DM PD_BUF Q RE SAE VDDHD VDDI VSSI WE Y[0] Y[1] 
+ Y[2] Y[3]
*.PININFO AWT2:I BIST2IO:I BLEQ:I BWEB:I BWEBM:I CKD:I D:I DM:I PD_BUF:I RE:I 
*.PININFO SAE:I WE:I Y[0]:I Y[1]:I Y[2]:I Y[3]:I Q:O BL[0]:B BL[1]:B BL[2]:B 
*.PININFO BL[3]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B VDDHD:B VDDI:B VSSI:B
MP10 VDDHD PD_BUF VDDI VDDI PCH L=65.0N W=2.5U M=2
XI213 WE VSSI VDDI NET65 S1AHSF400W40_AINV FN=1 WN=0.15U LN=0.06U FP=1 WP=0.15U LP=0.06U 
+ M=1
XI268 BLEQ VSSI VDDI BLEQI S1AHSF400W40_AINV FN=1 WN=0.25U LN=0.06U FP=1 WP=0.5U LP=0.06U 
+ M=1
XI214 NET65 VSSI VDDI WEI S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 WP=0.4U LP=0.06U 
+ M=1
XI215 NET53 VSSI VDDI REI S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 WP=0.4U LP=0.06U 
+ M=1
XI216 RE VSSI VDDI NET53 S1AHSF400W40_AINV FN=1 WN=0.15U LN=0.06U FP=1 WP=0.15U LP=0.06U 
+ M=1
XYPASS BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] BLEQI DL DLB REI 
+ VDDI VSSI WC WEI WT Y[0] Y[1] Y[2] Y[3] S1AHSF400W40_YPASS_M4_SB
XDOUT AWT2 AWTD BLEQI DL DLB PD_BUF Q SAE VDDHD VDDI VSSI S1AHSF400W40_DOUT_SB
XDIN AWTD BIST2IO BWEB BWEBM CKD D DM VDDHD VSSI WC WT S1AHSF400W40_DIN_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_IO_LD_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_IO_LD_SIM AWT2_LT AWT2_RT BIST2IO_LT BIST2IO_RT BLEQ_LT BLEQ_RT 
+ CKD_LT CKD_RT PD_BUF_LT PD_BUF_RT RE_LT RE_RT SAE_LT SAE_RT VDDHD VDDI VSSI 
+ WE_LT WE_RT YL_LT[0] YL_LT[1] YL_RT[0] YL_RT[1] Y_LT[0] Y_LT[1] Y_LT[2] 
+ Y_LT[3] Y_LT[4] Y_LT[5] Y_LT[6] Y_LT[7] Y_RT[0] Y_RT[1] Y_RT[2] Y_RT[3] 
+ Y_RT[4] Y_RT[5] Y_RT[6] Y_RT[7]
*.PININFO AWT2_LT:B AWT2_RT:B BIST2IO_LT:B BIST2IO_RT:B BLEQ_LT:B BLEQ_RT:B 
*.PININFO CKD_LT:B CKD_RT:B PD_BUF_LT:B PD_BUF_RT:B RE_LT:B RE_RT:B SAE_LT:B 
*.PININFO SAE_RT:B VDDHD:B VDDI:B VSSI:B WE_LT:B WE_RT:B YL_LT[0]:B YL_LT[1]:B 
*.PININFO YL_RT[0]:B YL_RT[1]:B Y_LT[0]:B Y_LT[1]:B Y_LT[2]:B Y_LT[3]:B 
*.PININFO Y_LT[4]:B Y_LT[5]:B Y_LT[6]:B Y_LT[7]:B Y_RT[0]:B Y_RT[1]:B 
*.PININFO Y_RT[2]:B Y_RT[3]:B Y_RT[4]:B Y_RT[5]:B Y_RT[6]:B Y_RT[7]:B
XI23 NET0160 NET0102 NET0146[0] NET0146[1] NET0146[2] NET0146[3] NET0146[4] 
+ NET0146[5] NET0146[6] NET0146[7] NET0146[8] NET0146[9] NET0146[10] 
+ NET0146[11] NET0146[12] NET0146[13] NET0146[14] NET0146[15] NET0134[0] 
+ NET0134[1] NET0134[2] NET0134[3] NET0134[4] NET0134[5] NET0134[6] NET0134[7] 
+ NET0134[8] NET0134[9] NET0134[10] NET0134[11] NET0134[12] NET0134[13] 
+ NET0134[14] NET0134[15] NET0148 NET0103 NET09 NET0157 NET0141 NET0149 NET090 
+ NET0139 NET06 NET0156 NET0130 NET0161 NET0143 NET0128 NET0165[0] NET0165[1] 
+ NET0165[2] NET0165[3] NET0165[4] NET0165[5] NET0165[6] NET0165[7] NET0145[0] 
+ NET0145[1] S1AHSF400W40_MIO_M16_SB
XI22 NET049 NET0131 NET0137[0] NET0137[1] NET0137[2] NET0137[3] NET0137[4] 
+ NET0137[5] NET0137[6] NET0137[7] NET0155[0] NET0155[1] NET0155[2] NET0155[3] 
+ NET0155[4] NET0155[5] NET0155[6] NET0155[7] NET0166 NET0152 NET0150 NET0158 
+ NET095 NET0136 NET0151 NET0101 NET0162 NET0106 NET0163 NET091 NET0153 
+ NET0132 NET048[0] NET048[1] NET048[2] NET048[3] NET048[4] NET048[5] 
+ NET048[6] NET048[7] S1AHSF400W40_MIO_M8_SB
XI21 NET0117 NET0112 NET0119[0] NET0119[1] NET0119[2] NET0119[3] NET0125[0] 
+ NET0125[1] NET0125[2] NET0125[3] NET0111 NET0116 NET0115 NET0120 NET0114 
+ NET0113 NET0122 NET0118 NET068 NET0124 NET0126 NET0121 NET0109 NET069 
+ NET070[0] NET070[1] NET070[2] NET070[3] S1AHSF400W40_MIO_M4_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    DIN_M16_BIST_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_DIN_M16_BIST_SB AWTD BIST BWEB BWEBM CKD D DM VDDHD VSSI WC[0] WC[1] 
+ WT[0] WT[1] YL[0] YL[1]
*.PININFO BIST:I BWEB:I BWEBM:I CKD:I D:I DM:I YL[0]:I YL[1]:I AWTD:O WC[0]:O 
*.PININFO WC[1]:O WT[0]:O WT[1]:O VDDHD:B VSSI:B
XI353 CKD1B VSSI VSSI VDDHD VDDHD CKD2 S1AHSF400W40_INV_BULK FN=1 WN=0.6U LN=0.06U FP=1 
+ WP=1.2U LP=0.06U M=1
XI354 CKD VSSI VSSI VDDHD VDDHD CKD1B S1AHSF400W40_INV_BULK FN=1 WN=0.4U LN=0.06U FP=1 
+ WP=0.8U LP=0.06U M=1
XI355 BIST1B VSSI VSSI VDDHD VDDHD BIST2 S1AHSF400W40_INV_BULK FN=1 WN=0.6U LN=0.06U FP=1 
+ WP=1.2U LP=0.06U M=1
XI356 BIST VSSI VSSI VDDHD VDDHD BIST1B S1AHSF400W40_INV_BULK FN=1 WN=0.4U LN=0.06U FP=1 
+ WP=0.8U LP=0.06U M=1
XI76 GWB YL[0] VSSI VDDHD NET249 S1AHSF400W40_ANAND FN2=1 WN2=0.5U LN2=0.06U FN1=1 
+ WN1=0.5U LN1=0.06U FP1=1 WP1=0.5U LP1=0.06U FP2=1 WP2=0.5U LP2=0.06U M=1
XI281 GW YL[1] VSSI VDDHD NET239 S1AHSF400W40_ANAND FN2=1 WN2=0.5U LN2=0.06U FN1=1 
+ WN1=0.5U LN1=0.06U FP1=1 WP1=0.5U LP1=0.06U FP2=1 WP2=0.5U LP2=0.06U M=1
XI280 GWB YL[1] VSSI VDDHD NET234 S1AHSF400W40_ANAND FN2=1 WN2=0.5U LN2=0.06U FN1=1 
+ WN1=0.5U LN1=0.06U FP1=1 WP1=0.5U LP1=0.06U FP2=1 WP2=0.5U LP2=0.06U M=1
XI279 GW YL[0] VSSI VDDHD NET244 S1AHSF400W40_ANAND FN2=1 WN2=0.5U LN2=0.06U FN1=1 
+ WN1=0.5U LN1=0.06U FP1=1 WP1=0.5U LP1=0.06U FP2=1 WP2=0.5U LP2=0.06U M=1
MM70 BXL CKD1B Z16 VDDHD PCH L=120.0N W=600N M=1
MM71 Z21 D VDDHD VDDHD PCH L=120.0N W=600N M=1
MM72 DXL DXB Z9 VDDHD PCH L=120.0N W=600N M=1
MM73 DXL CKD1B Z6 VDDHD PCH L=120.0N W=600N M=1
MM74 D_BIST BIST1B Z22 VDDHD PCH L=120.0N W=600N M=1
MM75 D_BIST BIST2 Z21 VDDHD PCH L=120.0N W=600N M=1
MM76 BXL BXB Z13 VDDHD PCH L=120.0N W=600N M=1
MP19 B_BIST BIST2 Z25 VDDHD PCH L=120.0N W=600N M=1
MM66 DXL3B_AND BXL1B VDDHD VDDHD PCH L=60N W=500N M=2
MP18 Z25 BWEB VDDHD VDDHD PCH L=120.0N W=600N M=1
MP16 B_BIST BIST1B Z26 VDDHD PCH L=120.0N W=600N M=1
MM61 DXL3B_AND DXL2 VDDHD VDDHD PCH L=60N W=500N M=2
MM62 VDDHD DXL1B Z6 VDDHD PCH L=120.0N W=600N M=1
MM63 Z22 DM VDDHD VDDHD PCH L=120.0N W=600N M=1
MP25 Z26 BWEBM VDDHD VDDHD PCH L=120.0N W=600N M=1
MP10 DXL2_AND CKD2 VDDHD VDDHD PCH L=60N W=500N M=2
MP1 DXL3B_AND CKD2 VDDHD VDDHD PCH L=60N W=500N M=2
MM64 DXL2_AND DXL1B VDDHD VDDHD PCH L=60N W=500N M=2
MM65 DXL2_AND BXL1B VDDHD VDDHD PCH L=60N W=500N M=2
MM67 VDDHD CKD2 Z9 VDDHD PCH L=120.0N W=600N M=1
MM68 VDDHD CKD2 Z13 VDDHD PCH L=120.0N W=600N M=1
MM69 VDDHD BXL1B Z16 VDDHD PCH L=120.0N W=600N M=1
MM55 DXL DXB Z11 VSSI NCH L=120.0N W=300N M=1
MM54 VSSI CKD1B Z11 VSSI NCH L=120.0N W=300N M=1
MN33 DXL3B_AND DXL2 Z2 VSSI NCH L=60N W=1U M=2
MM56 Z23 D VSSI VSSI NCH L=120.0N W=300N M=1
MM50 BXL CKD2 Z14 VSSI NCH L=120.0N W=300N M=1
MN7 Z1 BXL1B VSSI VSSI NCH L=60N W=1U M=2
MM57 D_BIST BIST1B Z23 VSSI NCH L=120.0N W=300N M=1
MN2 Z2 CKD2 Z1 VSSI NCH L=60N W=1U M=2
MN27 B_BIST BIST2 Z28 VSSI NCH L=120.0N W=300N M=1
MM58 VSSI DXL1B Z7 VSSI NCH L=120.0N W=300N M=1
MM59 VSSI CKD1B Z15 VSSI NCH L=120.0N W=300N M=1
MM60 BXL BXB Z15 VSSI NCH L=120.0N W=300N M=1
MN16 Z28 BWEBM VSSI VSSI NCH L=120.0N W=300N M=1
MN1 DXL2_AND DXL1B Z2 VSSI NCH L=60N W=1U M=2
MN19 B_BIST BIST1B Z27 VSSI NCH L=120.0N W=300N M=1
MN17 Z27 BWEB VSSI VSSI NCH L=120.0N W=300N M=1
MM51 DXL CKD2 Z7 VSSI NCH L=120.0N W=300N M=1
MM53 Z24 DM VSSI VSSI NCH L=120.0N W=300N M=1
MM52 D_BIST BIST2 Z24 VSSI NCH L=120.0N W=300N M=1
MM49 VSSI BXL1B Z14 VSSI NCH L=120.0N W=300N M=1
XI358 NET0499 VSSI VDDHD WT[0] S1AHSF400W40_AINV FN=6 WN=0.8U LN=0.06U FP=6 WP=0.3U 
+ LP=0.06U M=1
XI360 NET0491 VSSI VDDHD WT[1] S1AHSF400W40_AINV FN=6 WN=0.8U LN=0.06U FP=6 WP=0.3U 
+ LP=0.06U M=1
XI359 NET0511 VSSI VDDHD WC[0] S1AHSF400W40_AINV FN=6 WN=0.8U LN=0.06U FP=6 WP=0.3U 
+ LP=0.06U M=1
XI276 NET244 VSSI VDDHD NET0511 S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U 
+ LP=0.06U M=1
XI277 NET234 VSSI VDDHD NET0491 S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U 
+ LP=0.06U M=1
XI347 DXL2_AND VSSI VDDHD GWB S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U LP=0.06U 
+ M=1
XI361 NET0487 VSSI VDDHD WC[1] S1AHSF400W40_AINV FN=6 WN=0.8U LN=0.06U FP=6 WP=0.3U 
+ LP=0.06U M=1
XI349 BXL VSSI VDDHD BXL1B S1AHSF400W40_AINV FN=2 WN=0.3U LN=0.06U FP=2 WP=0.6U LP=0.06U 
+ M=1
XI350 B_BIST VSSI VDDHD NET0546 S1AHSF400W40_AINV FN=1 WN=0.3U LN=120N FP=1 WP=0.3U 
+ LP=120N M=1
XI351 DXL VSSI VDDHD DXL1B S1AHSF400W40_AINV FN=2 WN=0.3U LN=0.06U FP=2 WP=0.6U LP=0.06U 
+ M=1
XINV01 NET0570 VSSI VDDHD DXB S1AHSF400W40_AINV FN=1 WN=0.3U LN=120N FP=1 WP=0.3U LP=120N 
+ M=1
XI254 DXL3B_AND VSSI VDDHD GW S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U LP=0.06U 
+ M=1
XI352 NET0546 VSSI VDDHD BXB S1AHSF400W40_AINV FN=1 WN=0.3U LN=120N FP=1 WP=0.3U LP=120N 
+ M=1
XINV05 DXL1B VSSI VDDHD DXL2 S1AHSF400W40_AINV FN=2 WN=0.3U LN=0.06U FP=2 WP=0.6U 
+ LP=0.06U M=1
XINV00 D_BIST VSSI VDDHD NET0570 S1AHSF400W40_AINV FN=1 WN=0.3U LN=120N FP=1 WP=0.3U 
+ LP=120N M=1
XINV1 NET249 VSSI VDDHD NET0499 S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U 
+ LP=0.06U M=1
XI278 NET239 VSSI VDDHD NET0487 S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U 
+ LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MIO_M16_BIST_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MIO_M16_BIST_SB AWT2 BIST2IO BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] 
+ BL[7] BL[8] BL[9] BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BLB[0] BLB[1] 
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] 
+ BLB[12] BLB[13] BLB[14] BLB[15] BLEQ BWEB BWEBM CKD D DM PD_BUF Q RE SAE 
+ VDDHD VDDI VSSI WE Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7] YL[0] YL[1]
*.PININFO AWT2:I BIST2IO:I BLEQ:I BWEB:I BWEBM:I CKD:I D:I DM:I PD_BUF:I RE:I 
*.PININFO SAE:I WE:I Y[0]:I Y[1]:I Y[2]:I Y[3]:I Y[4]:I Y[5]:I Y[6]:I Y[7]:I 
*.PININFO YL[0]:I YL[1]:I Q:O BL[0]:B BL[1]:B BL[2]:B BL[3]:B BL[4]:B BL[5]:B 
*.PININFO BL[6]:B BL[7]:B BL[8]:B BL[9]:B BL[10]:B BL[11]:B BL[12]:B BL[13]:B 
*.PININFO BL[14]:B BL[15]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B BLB[4]:B 
*.PININFO BLB[5]:B BLB[6]:B BLB[7]:B BLB[8]:B BLB[9]:B BLB[10]:B BLB[11]:B 
*.PININFO BLB[12]:B BLB[13]:B BLB[14]:B BLB[15]:B VDDHD:B VDDI:B VSSI:B
XDIN AWTD BIST2IO BWEB BWEBM CKD D DM VDDHD VSSI WC[0] WC[1] WT[0] WT[1] YL[0] 
+ YL[1] S1AHSF400W40_DIN_M16_BIST_SB
MP10 VDDHD PD_BUF VDDI VDDI PCH L=65.0N W=2.5U M=2
XDOUT AWT2 AWTD BLEQI DL[0] DL[1] DLB[0] DLB[1] PD_BUF Q SAE VDDHD VDDI VSSI 
+ YL[0] YL[1] S1AHSF400W40_DOUT_M16_SB
XYPASS BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BLB[0] BLB[1] BLB[2] 
+ BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLEQI DL[0] DLB[0] REI VDDI VSSI WC[0] 
+ WEI WT[0] Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7] S1AHSF400W40_YPASS_M8_SB
XYPASS_1 BL[8] BL[9] BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BLB[8] BLB[9] 
+ BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15] BLEQI DL[1] DLB[1] REI VDDI 
+ VSSI WC[1] WEI WT[1] Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7] S1AHSF400W40_YPASS_M8_SB
XI184 BLEQ VSSI VDDI BLEQI S1AHSF400W40_AINV FN=4 WN=0.2U LN=0.06U FP=4 WP=0.4U LP=0.06U 
+ M=1
XI213 WE VSSI VDDI NET280 S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 WP=0.4U LP=0.06U 
+ M=1
XI214 NET280 VSSI VDDI WEI S1AHSF400W40_AINV FN=1 WN=0.4U LN=0.06U FP=1 WP=0.8U LP=0.06U 
+ M=1
XI215 NET268 VSSI VDDI REI S1AHSF400W40_AINV FN=1 WN=0.4U LN=0.06U FP=1 WP=0.8U LP=0.06U 
+ M=1
XI216 RE VSSI VDDI NET268 S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 WP=0.4U LP=0.06U 
+ M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    DIN_BIST_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_DIN_BIST_SB AWTD BIST BWEB BWEBM CKD D DM VDDHD VSSI WC WT
*.PININFO BIST:I BWEB:I BWEBM:I CKD:I D:I DM:I AWTD:O WC:O WT:O VDDHD:B VSSI:B
XI317 GWB VSSI VDDHD WT S1AHSF400W40_AINV FN=6 WN=0.8U LN=0.06U FP=6 WP=0.4U LP=0.06U M=1
XI319 BXL VSSI VDDHD BXL1B S1AHSF400W40_AINV FN=2 WN=0.3U LN=0.06U FP=2 WP=0.6U LP=0.06U 
+ M=1
XI315 B_BIST VSSI VDDHD NET297 S1AHSF400W40_AINV FN=1 WN=0.3U LN=120N FP=1 WP=0.3U 
+ LP=120N M=1
XI318 DXL VSSI VDDHD DXL1B S1AHSF400W40_AINV FN=2 WN=0.3U LN=0.06U FP=2 WP=0.6U LP=0.06U 
+ M=1
XINV01 NET329 VSSI VDDHD DXB S1AHSF400W40_AINV FN=1 WN=0.3U LN=120N FP=1 WP=0.3U LP=120N 
+ M=1
XI254 DXL3B_AND VSSI VDDHD GW S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U LP=0.06U 
+ M=1
XI267 DXL2_AND VSSI VDDHD GWB S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U LP=0.06U 
+ M=1
XI316 NET297 VSSI VDDHD BXB S1AHSF400W40_AINV FN=1 WN=0.3U LN=120N FP=1 WP=0.3U LP=120N 
+ M=1
XINV07 GW VSSI VDDHD WC S1AHSF400W40_AINV FN=6 WN=0.8U LN=0.06U FP=6 WP=0.4U LP=0.06U M=1
XINV05 DXL1B VSSI VDDHD DXL2 S1AHSF400W40_AINV FN=2 WN=0.3U LN=0.06U FP=2 WP=0.6U 
+ LP=0.06U M=1
XINV00 D_BIST VSSI VDDHD NET329 S1AHSF400W40_AINV FN=1 WN=0.3U LN=120N FP=1 WP=0.3U 
+ LP=120N M=1
MM44 VSSI BXL1B Z14 VSSI NCH L=120.0N W=300N M=1
MM45 BXL CKD2 Z14 VSSI NCH L=120.0N W=300N M=1
MN19 B_BIST BIST1B Z27 VSSI NCH L=120.0N W=300N M=1
MN7 Z1 BXL1B VSSI VSSI NCH L=60N W=1U M=2
MN17 Z27 BWEB VSSI VSSI NCH L=120.0N W=300N M=1
MN1 DXL2_AND DXL1B Z2 VSSI NCH L=60N W=1U M=2
MM35 DXL CKD2 Z7 VSSI NCH L=120.0N W=300N M=1
MN33 DXL3B_AND DXL2 Z2 VSSI NCH L=60N W=1U M=2
MM33 D_BIST BIST2 Z24 VSSI NCH L=120.0N W=300N M=1
MM32 Z24 DM VSSI VSSI NCH L=120.0N W=300N M=1
MM36 VSSI CKD1B Z11 VSSI NCH L=120.0N W=300N M=1
MM34 DXL DXB Z11 VSSI NCH L=120.0N W=300N M=1
MM31 Z23 D VSSI VSSI NCH L=120.0N W=300N M=1
MM30 D_BIST BIST1B Z23 VSSI NCH L=120.0N W=300N M=1
MN2 Z2 CKD2 Z1 VSSI NCH L=60N W=1U M=2
MN27 B_BIST BIST2 Z28 VSSI NCH L=120.0N W=300N M=1
MM37 VSSI DXL1B Z7 VSSI NCH L=120.0N W=300N M=1
MM43 VSSI CKD1B Z15 VSSI NCH L=120.0N W=300N M=1
MM42 BXL BXB Z15 VSSI NCH L=120.0N W=300N M=1
MN16 Z28 BWEBM VSSI VSSI NCH L=120.0N W=300N M=1
MP16 B_BIST BIST1B Z26 VDDHD PCH L=120.0N W=600N M=1
MM51 DXL3B_AND DXL2 VDDHD VDDHD PCH L=60N W=500N M=2
MM28 VDDHD DXL1B Z6 VDDHD PCH L=120.0N W=600N M=1
MM25 Z22 DM VDDHD VDDHD PCH L=120.0N W=600N M=1
MP25 Z26 BWEBM VDDHD VDDHD PCH L=120.0N W=600N M=1
MP10 DXL2_AND CKD2 VDDHD VDDHD PCH L=60N W=500N M=2
MP1 DXL3B_AND CKD2 VDDHD VDDHD PCH L=60N W=500N M=2
MM52 DXL2_AND DXL1B VDDHD VDDHD PCH L=60N W=500N M=2
MM53 DXL2_AND BXL1B VDDHD VDDHD PCH L=60N W=500N M=2
MM54 DXL3B_AND BXL1B VDDHD VDDHD PCH L=60N W=500N M=2
MM26 VDDHD CKD2 Z9 VDDHD PCH L=120.0N W=600N M=1
MM38 VDDHD CKD2 Z13 VDDHD PCH L=120.0N W=600N M=1
MM39 VDDHD BXL1B Z16 VDDHD PCH L=120.0N W=600N M=1
MM40 BXL CKD1B Z16 VDDHD PCH L=120.0N W=600N M=1
MM22 Z21 D VDDHD VDDHD PCH L=120.0N W=600N M=1
MM27 DXL DXB Z9 VDDHD PCH L=120.0N W=600N M=1
MM29 DXL CKD1B Z6 VDDHD PCH L=120.0N W=600N M=1
MM24 D_BIST BIST1B Z22 VDDHD PCH L=120.0N W=600N M=1
MM23 D_BIST BIST2 Z21 VDDHD PCH L=120.0N W=600N M=1
MM41 BXL BXB Z13 VDDHD PCH L=120.0N W=600N M=1
MP18 Z25 BWEB VDDHD VDDHD PCH L=120.0N W=600N M=1
MP19 B_BIST BIST2 Z25 VDDHD PCH L=120.0N W=600N M=1
XI324 CKD1B VSSI VSSI VDDHD VDDHD CKD2 S1AHSF400W40_INV_BULK FN=1 WN=0.6U LN=0.06U FP=1 
+ WP=1.2U LP=0.06U M=1
XI323 CKD VSSI VSSI VDDHD VDDHD CKD1B S1AHSF400W40_INV_BULK FN=1 WN=0.4U LN=0.06U FP=1 
+ WP=0.8U LP=0.06U M=1
XI326 BIST1B VSSI VSSI VDDHD VDDHD BIST2 S1AHSF400W40_INV_BULK FN=1 WN=0.6U LN=0.06U FP=1 
+ WP=1.2U LP=0.06U M=1
XI325 BIST VSSI VSSI VDDHD VDDHD BIST1B S1AHSF400W40_INV_BULK FN=1 WN=0.4U LN=0.06U FP=1 
+ WP=0.8U LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MIO_M8_BIST_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MIO_M8_BIST_SB AWT2 BIST2IO BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] 
+ BL[7] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLEQ BWEB 
+ BWEBM CKD D DM PD_BUF Q RE SAE VDDHD VDDI VSSI WE Y[0] Y[1] Y[2] Y[3] Y[4] 
+ Y[5] Y[6] Y[7] YL[0] YL[1]
*.PININFO AWT2:I BIST2IO:I BLEQ:I BWEB:I BWEBM:I CKD:I D:I DM:I PD_BUF:I RE:I 
*.PININFO SAE:I WE:I Y[0]:I Y[1]:I Y[2]:I Y[3]:I Y[4]:I Y[5]:I Y[6]:I Y[7]:I 
*.PININFO YL[0]:I YL[1]:I Q:O BL[0]:B BL[1]:B BL[2]:B BL[3]:B BL[4]:B BL[5]:B 
*.PININFO BL[6]:B BL[7]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B BLB[4]:B 
*.PININFO BLB[5]:B BLB[6]:B BLB[7]:B VDDHD:B VDDI:B VSSI:B
MP10 VDDHD PD_BUF VDDI VDDI PCH L=65.0N W=2.5U M=2
XDIN AWTD BIST2IO BWEB BWEBM CKD D DM VDDHD VSSI WC WT S1AHSF400W40_DIN_BIST_SB
XDOUT AWT2 AWTD BLEQI DL DLB PD_BUF Q SAE VDDHD VDDI VSSI S1AHSF400W40_DOUT_SB
XYPASS BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BLB[0] BLB[1] BLB[2] 
+ BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLEQI DL DLB REI VDDI VSSI WC WEI WT Y[0] 
+ Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7] S1AHSF400W40_YPASS_M8_SB
XI216 RE VSSI VDDI NET101 S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 WP=0.4U LP=0.06U 
+ M=1
XI215 NET101 VSSI VDDI REI S1AHSF400W40_AINV FN=1 WN=0.4U LN=0.06U FP=1 WP=0.8U LP=0.06U 
+ M=1
XI213 WE VSSI VDDI NET89 S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 WP=0.4U LP=0.06U M=1
XI184 BLEQ VSSI VDDI BLEQI S1AHSF400W40_AINV FN=2 WN=0.25U LN=0.06U FP=2 WP=0.5U LP=0.06U 
+ M=1
XI214 NET89 VSSI VDDI WEI S1AHSF400W40_AINV FN=1 WN=0.4U LN=0.06U FP=1 WP=0.8U LP=0.06U 
+ M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MIO_M4_BIST_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MIO_M4_BIST_SB AWT2 BIST2IO BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] 
+ BLB[2] BLB[3] BLEQ BWEB BWEBM CKD D DM PD_BUF Q RE SAE VDDHD VDDI VSSI WE 
+ Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7] YL[0] YL[1]
*.PININFO AWT2:I BIST2IO:I BLEQ:I BWEB:I BWEBM:I CKD:I D:I DM:I PD_BUF:I RE:I 
*.PININFO SAE:I WE:I Y[0]:I Y[1]:I Y[2]:I Y[3]:I Y[4]:I Y[5]:I Y[6]:I Y[7]:I 
*.PININFO YL[0]:I YL[1]:I Q:O BL[0]:B BL[1]:B BL[2]:B BL[3]:B BLB[0]:B 
*.PININFO BLB[1]:B BLB[2]:B BLB[3]:B VDDHD:B VDDI:B VSSI:B
MP10 VDDHD PD_BUF VDDI VDDI PCH L=65.0N W=2.5U M=2
XDIN AWTD BIST2IO BWEB BWEBM CKD D DM VDDHD VSSI WC WT S1AHSF400W40_DIN_BIST_SB
XI213 WE VSSI VDDI NET65 S1AHSF400W40_AINV FN=1 WN=0.15U LN=0.06U FP=1 WP=0.15U LP=0.06U 
+ M=1
XI268 BLEQ VSSI VDDI BLEQI S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 WP=0.48U LP=0.06U 
+ M=1
XI214 NET65 VSSI VDDI WEI S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 WP=0.4U LP=0.06U 
+ M=1
XI215 NET53 VSSI VDDI REI S1AHSF400W40_AINV FN=1 WN=0.2U LN=0.06U FP=1 WP=0.4U LP=0.06U 
+ M=1
XI216 RE VSSI VDDI NET53 S1AHSF400W40_AINV FN=1 WN=0.15U LN=0.06U FP=1 WP=0.15U LP=0.06U 
+ M=1
XYPASS BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] BLEQI DL DLB REI 
+ VDDI VSSI WC WEI WT Y[0] Y[1] Y[2] Y[3] S1AHSF400W40_YPASS_M4_SB
XDOUT AWT2 AWTD BLEQI DL DLB PD_BUF Q SAE VDDHD VDDI VSSI S1AHSF400W40_DOUT_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_IO_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_IO_SIM AWT2_LT AWT2_RT BIST2IO_LT BIST2IO_RT BL[0] BL[1] BL[2] 
+ BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10] BL[11] BL[12] BL[13] BL[14] 
+ BL[15] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] 
+ BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15] BLEQ_LT BLEQ_RT BWEB BWEBM 
+ CKD_LT CKD_RT D DM PD_BUF_LT PD_BUF_RT Q RE_LT RE_RT SAE_LT SAE_RT VDDHD 
+ VDDI VSSI WE_LT WE_RT YL_LT[0] YL_LT[1] YL_RT[0] YL_RT[1] Y_LT[0] Y_LT[1] 
+ Y_LT[2] Y_LT[3] Y_LT[4] Y_LT[5] Y_LT[6] Y_LT[7] Y_RT[0] Y_RT[1] Y_RT[2] 
+ Y_RT[3] Y_RT[4] Y_RT[5] Y_RT[6] Y_RT[7]
*.PININFO BWEB:I BWEBM:I D:I DM:I Q:O AWT2_LT:B AWT2_RT:B BIST2IO_LT:B 
*.PININFO BIST2IO_RT:B BL[0]:B BL[1]:B BL[2]:B BL[3]:B BL[4]:B BL[5]:B BL[6]:B 
*.PININFO BL[7]:B BL[8]:B BL[9]:B BL[10]:B BL[11]:B BL[12]:B BL[13]:B BL[14]:B 
*.PININFO BL[15]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B BLB[4]:B BLB[5]:B 
*.PININFO BLB[6]:B BLB[7]:B BLB[8]:B BLB[9]:B BLB[10]:B BLB[11]:B BLB[12]:B 
*.PININFO BLB[13]:B BLB[14]:B BLB[15]:B BLEQ_LT:B BLEQ_RT:B CKD_LT:B CKD_RT:B 
*.PININFO PD_BUF_LT:B PD_BUF_RT:B RE_LT:B RE_RT:B SAE_LT:B SAE_RT:B VDDHD:B 
*.PININFO VDDI:B VSSI:B WE_LT:B WE_RT:B YL_LT[0]:B YL_LT[1]:B YL_RT[0]:B 
*.PININFO YL_RT[1]:B Y_LT[0]:B Y_LT[1]:B Y_LT[2]:B Y_LT[3]:B Y_LT[4]:B 
*.PININFO Y_LT[5]:B Y_LT[6]:B Y_LT[7]:B Y_RT[0]:B Y_RT[1]:B Y_RT[2]:B 
*.PININFO Y_RT[3]:B Y_RT[4]:B Y_RT[5]:B Y_RT[6]:B Y_RT[7]:B
XI17 NET072 NET059 NET071[0] NET071[1] NET071[2] NET071[3] NET071[4] NET071[5] 
+ NET071[6] NET071[7] NET071[8] NET071[9] NET071[10] NET071[11] NET071[12] 
+ NET071[13] NET071[14] NET071[15] NET057[0] NET057[1] NET057[2] NET057[3] 
+ NET057[4] NET057[5] NET057[6] NET057[7] NET057[8] NET057[9] NET057[10] 
+ NET057[11] NET057[12] NET057[13] NET057[14] NET057[15] NET058 NET052 NET047 
+ NET016 NET061 NET060 NET030 NET020 NET068 NET073 NET025 NET069 NET056 NET08 
+ NET064[0] NET064[1] NET064[2] NET064[3] NET064[4] NET064[5] NET064[6] 
+ NET064[7] NET05[0] NET05[1] S1AHSF400W40_MIO_M16_BIST_SB
XI18 NET093 NET028 NET092[0] NET092[1] NET092[2] NET092[3] NET092[4] NET092[5] 
+ NET092[6] NET092[7] NET041[0] NET041[1] NET041[2] NET041[3] NET041[4] 
+ NET041[5] NET041[6] NET041[7] NET050 NET084 NET083 NET088 NET012 NET046 
+ NET091 NET086 NET089 NET033 NET049 NET090 NET042 NET087 NET085[0] NET085[1] 
+ NET085[2] NET085[3] NET085[4] NET085[5] NET085[6] NET085[7] NET044[0] 
+ NET044[1] S1AHSF400W40_MIO_M8_BIST_SB
XI19 NET0113 NET0101 NET040[0] NET040[1] NET040[2] NET040[3] NET018[0] 
+ NET018[1] NET018[2] NET018[3] NET043 NET053 NET029 NET027 NET02 NET021 
+ NET0111 NET039 NET0109 NET0114 NET0115 NET024 NET026 NET07 NET048[0] 
+ NET048[1] NET048[2] NET048[3] NET048[4] NET048[5] NET048[6] NET048[7] 
+ NET019[0] NET019[1] S1AHSF400W40_MIO_M4_BIST_SB
XI16 NET032 NET075 NET070[0] NET070[1] NET070[2] NET070[3] NET070[4] NET070[5] 
+ NET070[6] NET070[7] NET070[8] NET070[9] NET070[10] NET070[11] NET070[12] 
+ NET070[13] NET070[14] NET070[15] NET0117[0] NET0117[1] NET0117[2] NET0117[3] 
+ NET0117[4] NET0117[5] NET0117[6] NET0117[7] NET0117[8] NET0117[9] 
+ NET0117[10] NET0117[11] NET0117[12] NET0117[13] NET0117[14] NET0117[15] 
+ NET074 NET079 NET078 NET082 NET077 NET076 NET0124 NET080 NET0125 NET0122 
+ NET063 NET0123 NET0108 NET081 NET0120[0] NET0120[1] NET0120[2] NET0120[3] 
+ NET0120[4] NET0120[5] NET0120[6] NET0120[7] NET015[0] NET015[1] S1AHSF400W40_MIO_M16_SB
XI15 NET010 NET0126 NET0110[0] NET0110[1] NET0110[2] NET0110[3] NET0110[4] 
+ NET0110[5] NET0110[6] NET0110[7] NET022[0] NET022[1] NET022[2] NET022[3] 
+ NET022[4] NET022[5] NET022[6] NET022[7] NET095 NET0121 NET01 NET031 NET062 
+ NET0119 NET051 NET045 NET0112 NET0106 NET0107 NET036 NET013 NET0127 NET03[0] 
+ NET03[1] NET03[2] NET03[3] NET03[4] NET03[5] NET03[6] NET03[7] S1AHSF400W40_MIO_M8_SB
XI14 NET066 NET065 NET097[0] NET097[1] NET097[2] NET097[3] NET098[0] NET098[1] 
+ NET098[2] NET098[3] NET0100 NET094 NET096 NET035 NET0103 NET034 NET067 
+ NET037 NET011 NET099 NET0104 NET0102 NET038 NET023 NET0105[0] NET0105[1] 
+ NET0105[2] NET0105[3] S1AHSF400W40_MIO_M4_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    WEBBUF_BIST_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_WEBBUF_BIST_SB BIST1B BIST2 CKC CKT VDDHD VSSI WEB WEBM WEBXL WEBXL1B
*.PININFO BIST1B:I BIST2:I CKC:I CKT:I WEB:I WEBM:I WEBXL:O WEBXL1B:O VDDHD:B 
*.PININFO VSSI:B
MM14 WEBX BIST1B N3 VDDHD PCH L=60N W=600N M=1
MM15 N3 WEBM VDDHD VDDHD PCH L=60N W=600N M=1
MM20 WEBXL CKC NET0115 VDDHD PCH L=60N W=300N M=1
MM21 NET0115 WEBXL1B VDDHD VDDHD PCH L=60N W=300N M=1
MM16 N5 CKT VDDHD VDDHD PCH L=60N W=1U M=2
MM6 WEBXL WEBX N5 VDDHD PCH L=60N W=1U M=2
MM8 WEBX BIST2 N1 VDDHD PCH L=60N W=600N M=1
MM10 N1 WEB VDDHD VDDHD PCH L=60N W=600N M=1
MM9 WEBX BIST1B N2 VSSI NCH L=60N W=300N M=1
MM11 N4 WEBM VSSI VSSI NCH L=60N W=300N M=1
MM13 WEBX BIST2 N4 VSSI NCH L=60N W=300N M=1
MM0 WEBXL WEBX N7 VSSI NCH L=60N W=1U M=2
MM19 WEBXL CKT NET076 VSSI NCH L=60N W=200N M=1
MM18 NET076 WEBXL1B VSSI VSSI NCH L=60N W=200N M=1
MM12 N2 WEB VSSI VSSI NCH L=60N W=300N M=1
MM17 N7 CKC VSSI VSSI NCH L=60N W=1U M=2
XI25 WEBXL VSSI VDDHD WEBXL1B S1AHSF400W40_AINV FN=2 WN=0.55U LN=0.06U FP=2 WP=1U 
+ LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    VHILO_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_VHILO_SB VDDHD VHI VLO VSSI
*.PININFO VHI:O VLO:O VDDHD:B VSSI:B
MP0 Z2 Z2 VDDHD VDDHD PCH L=60N W=600N M=1
MP2 VHI Z1 VDDHD VDDHD PCH L=60N W=600N M=10
MP7 Z2 Z1 VDDHD VDDHD PCH L=60N W=600N M=1
MN3 VSSI Z2 Z1 VSSI NCH L=60N W=600N M=1
MN1 VSSI Z2 VLO VSSI NCH L=60N W=1.2U M=10
MN0 VSSI Z1 Z1 VSSI NCH L=60N W=600N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65_LOGIC
* CELL NAME:    ANAND3
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ANAND3 A B C G V Y
*.PININFO A:I B:I C:I G:I V:I Y:O
M1 Y C V V PCH L=LP3 W=WP3 M=1*FP3
M4 Y B V V PCH L=LP2 W=WP2 M=1*FP2
M6 Y A V V PCH L=LP1 W=WP1 M=1*FP1
M8 NET14 A G G NCH L=LN1 W=WN1 M=1*FN1
M10 NET17 B NET14 G NCH L=LN2 W=WN2 M=1*FN2
M12 Y C NET17 G NCH L=LN3 W=WN3 M=1*FN3
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CKG_882_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CKG_882_SB CKP CLK EN RSC RSTCK TM VDDHD VSSI
*.PININFO CLK:I EN:I RSTCK:I TM:I CKP:O RSC:O VDDHD:B VSSI:B
XINV0 Z17 VSSI VDDHD RSCI S1AHSF400W40_AINV FN=3 WN=0.35U LN=0.06U FP=3 WP=0.7U LP=0.06U 
+ M=1
XI50 RSTCK CKP VSSI VDDHD RSC S1AHSF400W40_ANAND FN2=1 WN2=2U LN2=0.06U FN1=1 WN1=2U 
+ LN1=0.06U FP1=1 WP1=2U LP1=0.06U FP2=1 WP2=2U LP2=0.06U M=1
XNAND4 CKPC Z19 VSSI VDDHD CKP S1AHSF400W40_ANAND FN2=4 WN2=0.75U LN2=0.06U FN1=4 
+ WN1=0.75U LN1=0.06U FP1=4 WP1=3U LP1=0.06U FP2=4 WP2=1.5U LP2=0.06U M=1
XNAND5 CKP RSCI VSSI VDDHD Z19 S1AHSF400W40_ANAND FN2=1 WN2=0.54U LN2=0.06U FN1=1 
+ WN1=0.54U LN1=0.06U FP1=1 WP1=0.75U LP1=0.06U FP2=1 WP2=0.75U LP2=0.06U M=1
XNAND3 Z16 Z14 VSSI VDDHD Z17 S1AHSF400W40_ANAND FN2=1 WN2=0.54U LN2=0.06U FN1=1 
+ WN1=0.54U LN1=0.06U FP1=1 WP1=0.54U LP1=0.06U FP2=1 WP2=0.54U LP2=0.06U M=1
XI49 Z17 CLK VSSI VDDHD Z14 S1AHSF400W40_ANAND FN2=1 WN2=0.4U LN2=0.06U FN1=1 WN1=0.4U 
+ LN1=0.06U FP1=1 WP1=0.4U LP1=0.06U FP2=1 WP2=0.4U LP2=0.06U M=1
XNAND0 TM CLK VSSI VDDHD Z15 S1AHSF400W40_ANAND FN2=1 WN2=0.4U LN2=0.06U FN1=1 WN1=0.4U 
+ LN1=0.06U FP1=1 WP1=0.4U LP1=0.06U FP2=1 WP2=0.4U LP2=0.06U M=1
XNAND12 CLK RSCI EN VSSI VDDHD CKPC S1AHSF400W40_ANAND3 FN3=1 WN3=2U LN3=0.06U FN2=1 
+ WN2=2U LN2=0.06U FN1=1 WN1=2U LN1=0.06U FP1=1 WP1=1U LP1=0.06U FP2=1 WP2=1U 
+ LP2=0.06U FP3=1 WP3=1U LP3=0.06U M=1
XI53 RSTCK CKP Z15 VSSI VDDHD Z16 S1AHSF400W40_ANAND3 FN3=1 WN3=0.9U LN3=0.06U FN2=1 
+ WN2=0.9U LN2=0.06U FN1=1 WN1=0.9U LN1=0.06U FP1=1 WP1=0.6U LP1=0.06U FP2=1 
+ WP2=0.6U LP2=0.06U FP3=1 WP3=0.6U LP3=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65_LOGIC
* CELL NAME:    ANOR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ANOR A B G V Y
*.PININFO A:I B:I G:I V:I Y:O
M1 Y B NET021 V PCH L=LP2 W=WP2 M=1*FP2
M3 NET021 A V V PCH L=LP1 W=WP1 M=1*FP1
M5 Y A G G NCH L=LN1 W=WN1 M=1*FN1
M7 Y B G G NCH L=LN2 W=WN2 M=1*FN2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    RESETD_TSEL
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_RESETD_TSEL CKP V[0] V[1] VDDHD VSSI TD_01_11 TD_10
*.PININFO CKP:I V[0]:I V[1]:I TD_01_11:O TD_10:O VDDHD:B VSSI:B
XI21 CKP VSSI VDDHD Z3 S1AHSF400W40_AINV FN=1 WN=0.3U LN=60N FP=1 WP=0.6U LP=60N M=1
XI78 Z4 VSSI VDDHD Z5 S1AHSF400W40_AINV FN=1 WN=0.3U LN=60N FP=1 WP=0.6U LP=60N M=1
XI77 Z3 VSSI VDDHD Z4 S1AHSF400W40_AINV FN=1 WN=0.3U LN=60N FP=1 WP=0.6U LP=60N M=1
XND0 CKP TD_10 VSSI VDDHD Z0 S1AHSF400W40_ANAND FN2=1 WN2=0.6U LN2=0.06U FN1=1 WN1=0.6U 
+ LN1=0.06U FP1=1 WP1=0.6U LP1=0.06U FP2=1 WP2=0.6U LP2=0.06U M=1
XI76 Z0 V[0] VSSI VDDHD TD_01_11 S1AHSF400W40_ANAND FN2=1 WN2=0.6U LN2=0.06U FN1=1 
+ WN1=0.6U LN1=0.06U FP1=1 WP1=0.6U LP1=0.06U FP2=1 WP2=0.6U LP2=0.06U M=1
XI79 Z5 V[1] VSSI VDDHD TD_10 S1AHSF400W40_ANAND FN2=1 WN2=0.6U LN2=0.06U FN1=1 WN1=0.6U 
+ LN1=0.06U FP1=1 WP1=0.6U LP1=0.06U FP2=1 WP2=0.6U LP2=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    RESETD_882_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_RESETD_882_SB BLTRKWLDRV CK2 CKP CKPD CKPDCLK DEC_X2[0] DEC_X2[1] 
+ IOSAEB RSTCK TK TRKBL VDDHD VSSI WEBXL WLP_SAE WLP_SAE_TK PTSEL RV[0] RV[1] 
+ WV[0] WV[1] WV[2]
*.PININFO CK2:I CKP:I DEC_X2[0]:I DEC_X2[1]:I WEBXL:I PTSEL:I RV[0]:I RV[1]:I 
*.PININFO WV[0]:I WV[1]:I WV[2]:I BLTRKWLDRV:O CKPD:O CKPDCLK:O IOSAEB:O 
*.PININFO RSTCK:O WLP_SAE:O TK:B TRKBL:B VDDHD:B VSSI:B WLP_SAE_TK:B
XI28 DEC_X2[0] DEC_X2[1] VSSI VDDHD DEC_NOR1B S1AHSF400W40_ANOR FN2=1 WN2=0.3U LN2=0.06U 
+ FN1=1 WN1=0.3U LN1=0.06U FP1=1 WP1=0.6U LP1=0.06U FP2=1 WP2=0.6U LP2=0.06U 
+ M=1
XTSEL_WT BLTRKWLDRV WV[0] WV[1] VDDHD VSSI NET118 NET115 S1AHSF400W40_RESETD_TSEL
XTSEL_RT CKP RV[0] RV[1] VDDHD VSSI RTD_01_11 RTD_10 S1AHSF400W40_RESETD_TSEL
XI673 DEC_NOR1B VSSI VDDHD NET0168 S1AHSF400W40_AINV FN=1 WN=0.4U LN=60N FP=1 WP=0.8U 
+ LP=60N M=1
XI537 RTKB2 VSSI VDDHD BLTRKWLDRV S1AHSF400W40_AINV FN=12 WN=0.5U LN=60N FP=6 WP=2U 
+ LP=60N M=1
XI668 SHORT_D1 VSSI VDDHD NET0145 S1AHSF400W40_AINV FN=1 WN=0.4U LN=60N FP=1 WP=0.8U 
+ LP=60N M=1
XI653 SAE_FIRE2 VSSI VDDHD WLP_SAE S1AHSF400W40_AINV FN=12 WN=0.5U LN=60N FP=6 WP=2U 
+ LP=60N M=1
XI594 Z1 VSSI VDDHD CKPD S1AHSF400W40_AINV FN=8 WN=0.5U LN=0.06U FP=4 WP=2U LP=0.06U M=1
XI593 CKP VSSI VDDHD Z1 S1AHSF400W40_AINV FN=1 WN=1U LN=0.06U FP=1 WP=2U LP=0.06U M=1
XI541 RTKB VSSI VDDHD RTKB1B S1AHSF400W40_AINV FN=2 WN=0.4U LN=60N FP=2 WP=0.8U LP=60N M=1
XI574 VDDHD VSSI VDDHD TRKBL1B S1AHSF400W40_AINV FN=3 WN=0.35U LN=90N FP=3 WP=0.7U LP=90N 
+ M=1
XI540 RTKB1B VSSI VDDHD RTKB2 S1AHSF400W40_AINV FN=6 WN=0.4U LN=60N FP=6 WP=0.8U LP=60N 
+ M=1
XI661 TRKBL1B VSSI VDDHD NET0184 S1AHSF400W40_AINV FN=2 WN=0.25U LN=60N FP=2 WP=0.5U 
+ LP=60N M=1
XI669 NET0145 VSSI VDDHD SHORT_D2 S1AHSF400W40_AINV FN=1 WN=0.4U LN=60N FP=1 WP=0.8U 
+ LP=60N M=1
XI666 SHORT_D2 TRKBL VSSI VDDHD NET168 S1AHSF400W40_ANAND FN2=2 WN2=0.5U LN2=90N FN1=2 
+ WN1=0.5U LN1=60N FP1=2 WP1=0.5U LP1=60N FP2=2 WP2=0.5U LP2=90N M=1
XI658 WV[2] RTKB1B VSSI VDDHD SHORT_D1 S1AHSF400W40_ANAND FN2=1 WN2=0.6U LN2=60N FN1=1 
+ WN1=0.6U LN1=60N FP1=1 WP1=0.6U LP1=60N FP2=1 WP2=0.6U LP2=60N M=1
XI654 SHORT_D1 NET0187 VSSI VDDHD RSTCK S1AHSF400W40_ANAND FN2=2 WN2=0.75U LN2=60N FN1=2 
+ WN1=0.75U LN1=60N FP1=2 WP1=0.75U LP1=60N FP2=2 WP2=0.75U LP2=60N M=1
XI667 WEBXL BLTRKWLDRV NET168 VSSI VDDHD SAE_FIRE2 S1AHSF400W40_ANAND3 FN3=1 WN3=3U 
+ LN3=60N FN2=1 WN2=3U LN2=60N FN1=1 WN1=3U LN1=60N FP1=1 WP1=3U LP1=60N FP2=1 
+ WP2=3U LP2=60N FP3=1 WP3=3U LP3=60N M=1
XI664 BLTRKWLDRV NET118 NET115 VSSI VDDHD NET0187 S1AHSF400W40_ANAND3 FN3=1 WN3=0.6U 
+ LN3=60N FN2=1 WN2=0.6U LN2=60N FN1=1 WN1=0.6U LN1=60N FP1=1 WP1=0.6U LP1=60N 
+ FP2=1 WP2=0.6U LP2=60N FP3=1 WP3=0.6U LP3=60N M=1
XI584 CKP RTD_01_11 RTD_10 VSSI VDDHD RTKB S1AHSF400W40_ANAND3 FN3=2 WN3=0.6U LN3=60N 
+ FN2=2 WN2=0.6U LN2=60N FN1=2 WN1=0.6U LN1=60N FP1=2 WP1=0.4U LP1=60N FP2=2 
+ WP2=0.4U LP2=60N FP3=2 WP3=0.4U LP3=60N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    BISTD_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BISTD_SB BIST BIST1B BIST2 BIST2IO VDDHD VSSI
*.PININFO BIST:I BIST1B:O BIST2:O BIST2IO:O VDDHD:B VSSI:B
XINV2 BIST1B_2 VSSI VDDHD BIST2 S1AHSF400W40_AINV FN=3 WN=1U LN=0.06U FP=3 WP=2U LP=0.06U 
+ M=1
XINV1 BIST VSSI VDDHD BIST1B_2 S1AHSF400W40_AINV FN=1 WN=1U LN=0.06U FP=1 WP=2U LP=0.06U 
+ M=1
XINV3 BIST1B_2 VSSI VDDHD BIST2IO S1AHSF400W40_AINV FN=6 WN=1U LN=0.06U FP=6 WP=2U 
+ LP=0.06U M=1
XI21 BIST VSSI VDDHD BIST1B S1AHSF400W40_AINV FN=3 WN=1U LN=0.06U FP=3 WP=2U LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    PDBUF_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_PDBUF_SB PD PDBUF VDDI VSSI
*.PININFO PD:I PDBUF:O VDDI:B VSSI:B
XINV0 PD VSSI VDDI NET37 S1AHSF400W40_AINV FN=2 WN=1U LN=0.06U FP=2 WP=1.5U LP=0.06U M=1
XINV2 NET37 VSSI VDDI PDBUF S1AHSF400W40_AINV FN=8 WN=1U LN=0.06U FP=8 WP=1.5U LP=0.06U 
+ M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    COTH_BIST_882_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_COTH_BIST_882_SB AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B 
+ CK2 CKP CKPD CLK DEC_X2[0] DEC_X2[1] EN PD PD_BUF PTSEL RSC RTSEL[0] 
+ RTSEL[1] TK TM TRKBL VDDHD VDDI VHI VLO VSSI WEB WEBM WEBXL WEBXL1B WLP_SAE 
+ WLP_SAEB WLP_SAE_TK WTSEL[0] WTSEL[1] WTSEL[2]
*.PININFO AWT:I BIST:I CK1B:I CK2:I CLK:I DEC_X2[0]:I DEC_X2[1]:I EN:I PD:I 
*.PININFO PTSEL:I RTSEL[0]:I RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I 
*.PININFO WTSEL[1]:I WTSEL[2]:I AWT2:O BIST1B:O BIST2:O BIST2IO:O BLTRKWLDRV:O 
*.PININFO CKP:O CKPD:O PD_BUF:O RSC:O VHI:O VLO:O WEBXL:O WEBXL1B:O WLP_SAE:O 
*.PININFO WLP_SAEB:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE_TK:B
MP1 VDDHD PD VDDI VDDI PCH L=60N W=3U M=22
MP0 VDDHD PD VDDI VDDI PCH L=60N W=3.8U M=29
XWEBBUF BIST1B BIST2 CK1B CK2 VDDHD VSSI WEB WEBM WEBXL WEBXL1B 
+ S1AHSF400W40_WEBBUF_BIST_SB
XVHILO_SB VDDHD VHI VLO VSSI S1AHSF400W40_VHILO_SB
XCKG CKP CLK EN RSC RSTCK TM VDDHD VSSI S1AHSF400W40_CKG_882_SB
XRESETD BLTRKWLDRV CK2 CKP CKPD CKPDCLK DEC_X2[0] DEC_X2[1] WLP_SAEB RSTCK TK 
+ TRKBL VDDHD VSSI WEBXL WLP_SAE WLP_SAE_TK PTSEL RTSEL[0] RTSEL[1] WTSEL[0] 
+ WTSEL[1] WTSEL[2] S1AHSF400W40_RESETD_882_SB
XBISTD_SB BIST BIST1B BIST2 BIST2IO VDDHD VSSI S1AHSF400W40_BISTD_SB
XPDBUF_SB PD PD_BUF VDDI VSSI S1AHSF400W40_PDBUF_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    DECB4_882_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_DECB4_882_SB IN0A IN0B IN1A IN1B IN2 PD PREDEC0 PREDEC1 PREDEC2 
+ PREDEC3 VDDHD VSSI
*.PININFO IN0A:I IN0B:I IN1A:I IN1B:I IN2:I PD:I PREDEC0:O PREDEC1:O PREDEC2:O 
*.PININFO PREDEC3:O VDDHD:B VSSI:B
MM6 PREDEC0 PD VSSI VSSI NCH L=60N W=300N M=1
MM11 PREDEC3 PD VSSI VSSI NCH L=60N W=300N M=1
MM10 PREDEC2 PD VSSI VSSI NCH L=60N W=300N M=1
MM3 NET137 IN2 VSSI VSSI NCH L=60N W=600N M=4
MM9 PREDEC1 PD VSSI VSSI NCH L=60N W=300N M=1
MM0 N1 IN0A N2 VSSI NCH L=60N W=600N M=1
MM7 N3 IN0B N2 VSSI NCH L=60N W=600N M=1
MM8 N2 IN1A NET137 VSSI NCH L=60N W=600N M=2
MM21 N4 IN0A N5 VSSI NCH L=60N W=600N M=1
MM20 N6 IN0B N5 VSSI NCH L=60N W=600N M=1
MM19 N5 IN1B NET137 VSSI NCH L=60N W=600N M=2
MM1 N1 IN0A VDDHD VDDHD PCH L=60N W=600N M=1
MM2 N1 IN1A VDDHD VDDHD PCH L=60N W=600N M=1
MM4 N3 IN0B VDDHD VDDHD PCH L=60N W=600N M=1
MM5 N3 IN1A VDDHD VDDHD PCH L=60N W=600N M=1
MM25 N1 IN2 VDDHD VDDHD PCH L=60N W=600N M=2
MM24 N3 IN2 VDDHD VDDHD PCH L=60N W=600N M=2
MM23 N6 IN2 VDDHD VDDHD PCH L=60N W=600N M=2
MM22 N4 IN2 VDDHD VDDHD PCH L=60N W=600N M=2
MM18 N4 IN0A VDDHD VDDHD PCH L=60N W=600N M=1
MM17 N4 IN1B VDDHD VDDHD PCH L=60N W=600N M=1
MM16 N6 IN0B VDDHD VDDHD PCH L=60N W=600N M=1
MM15 N6 IN1B VDDHD VDDHD PCH L=60N W=600N M=1
XINV0 N1 VSSI VDDHD PREDEC0 S1AHSF400W40_AINV FN=4 WN=0.7U LN=0.06U FP=4 WP=1.4U LP=0.06U 
+ M=1
XINV1 N3 VSSI VDDHD PREDEC1 S1AHSF400W40_AINV FN=4 WN=0.7U LN=0.06U FP=4 WP=1.4U LP=0.06U 
+ M=1
XINV2 N4 VSSI VDDHD PREDEC2 S1AHSF400W40_AINV FN=4 WN=0.7U LN=0.06U FP=4 WP=1.4U LP=0.06U 
+ M=1
XINV3 N6 VSSI VDDHD PREDEC3 S1AHSF400W40_AINV FN=4 WN=0.7U LN=0.06U FP=4 WP=1.4U LP=0.06U 
+ M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    ENBUFB_BIST_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ENBUFB_BIST_SB BIST1B BIST2 CEB CEBM CK1B CK2 CKP CLK CLK_ENV EN ENC 
+ RSC VDDHD VSSI
*.PININFO BIST1B:I BIST2:I CEB:I CEBM:I CK1B:I CK2:I CKP:I CLK:I RSC:I 
*.PININFO CLK_ENV:O EN:O ENC:O VDDHD:B VSSI:B
MM21 VDDHD EN ENC VDDHD PCH L=60N W=700N M=3
MM14 CEBX BIST1B NET0126 VDDHD PCH L=60N W=500N M=1
MM6 VDDHD CKP CLK_ENV VDDHD PCH L=60N W=750.0N M=4
MM1 CEBXL CK1B NET0158 VDDHD PCH L=60N W=500N M=1
MM16 CEBXL CEBX N5 VDDHD PCH L=60N W=1U M=2
MM7 CEBXL RSC VDDHD VDDHD PCH L=60N W=700N M=2
MM15 NET0126 CEBM VDDHD VDDHD PCH L=60N W=500N M=1
MM2 NET0158 EN VDDHD VDDHD PCH L=60N W=500N M=1
MM19 N5 CK2 VDDHD VDDHD PCH L=60N W=1U M=2
MM8 CEBX BIST2 NET0134 VDDHD PCH L=60N W=500N M=1
MM10 NET0134 CEB VDDHD VDDHD PCH L=60N W=500N M=1
MM22 ENC CLK NET0155 VSSI NCH L=60N W=3.2U M=5
MM23 ENC CKP NET0155 VSSI NCH L=60N W=3.2U M=1
MM0 NET0155 EN VSSI VSSI NCH L=60N W=3.2U M=5
MM18 N7 CK1B NET0187 VSSI NCH L=60N W=1U M=1
MM11 NET0195 CEBM VSSI VSSI NCH L=60N W=500N M=1
MM17 CEBXL CEBX N7 VSSI NCH L=60N W=1U M=1
MM20 NET0187 RSC VSSI VSSI NCH L=60N W=1U M=2
MM3 CEBXL CK2 NET0179 VSSI NCH L=60N W=500N M=1
MM12 NET0163 CEB VSSI VSSI NCH L=60N W=500N M=1
MM4 NET0179 EN NET0171 VSSI NCH L=60N W=500N M=1
MM9 CEBX BIST1B NET0163 VSSI NCH L=60N W=500N M=1
MM5 NET0171 RSC VSSI VSSI NCH L=60N W=1U M=1
MM13 CEBX BIST2 NET0195 VSSI NCH L=60N W=500N M=1
XI141 CEBXL VSSI VDDHD EN S1AHSF400W40_AINV FN=3 WN=1U LN=0.06U FP=3 WP=2U LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    ABUF_BIST_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ABUF_BIST_SB A AM AX1B AX1BL AX1BL1B BIST1B BIST2 CK1B CK2 VDDHD VSSI
*.PININFO A:I AM:I BIST1B:I BIST2:I CK1B:I CK2:I AX1B:O AX1BL:O AX1BL1B:O 
*.PININFO VDDHD:B VSSI:B
MM26 AX1BL CK1B NET94 VDDHD PCH L=60N W=300N M=1
MM24 AX BIST1B NET095 VDDHD PCH L=60N W=600N M=1
MM28 N5 CK2 VDDHD VDDHD PCH L=60N W=1U M=2
MM30 AX BIST2 N1 VDDHD PCH L=60N W=600N M=1
MM25 NET095 AM VDDHD VDDHD PCH L=60N W=600N M=1
MM27 NET94 AX1BL1B VDDHD VDDHD PCH L=60N W=300N M=1
MM29 AX1BL AX1B N5 VDDHD PCH L=60N W=1U M=2
MM31 N1 A VDDHD VDDHD PCH L=60N W=600N M=1
MM20 AX1BL CK2 NET111 VSSI NCH L=60N W=200N M=1
MM16 AX BIST1B N3 VSSI NCH L=60N W=300N M=1
MM23 N7 CK1B VSSI VSSI NCH L=60N W=1U M=2
MM19 AX1BL AX1B N7 VSSI NCH L=60N W=1U M=2
MM22 N3 A VSSI VSSI NCH L=60N W=300N M=1
MM17 NET0140 AM VSSI VSSI NCH L=60N W=300N M=1
MM18 AX BIST2 NET0140 VSSI NCH L=60N W=300N M=1
MM21 NET111 AX1BL1B VSSI VSSI NCH L=60N W=200N M=1
XI25 AX1BL VSSI VDDHD AX1BL1B S1AHSF400W40_AINV FN=1 WN=0.55U LN=0.06U FP=1 WP=1.0U 
+ LP=0.06U M=1
XI39 AX VSSI VDDHD AX1B S1AHSF400W40_AINV FN=4 WN=0.15U LN=0.06U FP=4 WP=0.25U LP=0.06U 
+ M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    DECB1_X_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_DECB1_X_SB CKP CLK DEC EN ENC PD PREDEC VDDHD VSSI
*.PININFO CKP:I CLK:I EN:I ENC:I PD:I PREDEC:I DEC:O VDDHD:B VSSI:B
MM0 NT1 PREDEC VDDHD VDDHD PCH L=60N W=1.25U M=2
MP0 DEC NT1 VDDHD VDDHD PCH L=60N W=2.5U M=4
MM1 NT1 PREDEC VSSI VSSI NCH L=60N W=625.00N M=2
MM5 DEC PD VSSI VSSI NCH L=60N W=300N M=1
MN0 DEC NT1 VSSI VSSI NCH L=60N W=2.5U M=2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    DECB1_BLEQ_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_DECB1_BLEQ_SB BLEQ CLK CLK_ENV ENC EN_DCLK PD VDDHD VDDI VSSI
*.PININFO CLK:I CLK_ENV:I ENC:I EN_DCLK:I PD:I BLEQ:O VDDHD:B VDDI:B VSSI:B
MP5 VDDHD EN_DCLK ENC VDDHD PCH L=60N W=800N M=4
MM2 CLK_ENV CLK ENC VDDHD PCH L=60N W=250.0N M=8
MP1 BLEQ ENC VDDHD VDDHD PCH L=60N W=2.5U M=8
MM5 BLEQ PD VSSI VSSI NCH L=60N W=300N M=2
MN1 BLEQ ENC VSSI VSSI NCH L=60N W=1.25U M=8
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    DECB4_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_DECB4_SB IN0A IN0B IN1A IN1B IN2 PREDEC0 PREDEC1 PREDEC2 PREDEC3 VDDHD 
+ VSSI
*.PININFO IN0A:I IN0B:I IN1A:I IN1B:I IN2:I PREDEC0:O PREDEC1:O PREDEC2:O 
*.PININFO PREDEC3:O VDDHD:B VSSI:B
MM3 NET137 IN2 VSSI VSSI NCH L=60N W=600N M=4
MM0 N1 IN0A N2 VSSI NCH L=60N W=600N M=1
MM7 N3 IN0B N2 VSSI NCH L=60N W=600N M=1
MM8 N2 IN1A NET137 VSSI NCH L=60N W=600N M=2
MM21 N4 IN0A N5 VSSI NCH L=60N W=600N M=1
MM20 N6 IN0B N5 VSSI NCH L=60N W=600N M=1
MM19 N5 IN1B NET137 VSSI NCH L=60N W=600N M=2
MM1 N1 IN0A VDDHD VDDHD PCH L=60N W=600N M=1
MM2 N1 IN1A VDDHD VDDHD PCH L=60N W=600N M=1
MM4 N3 IN0B VDDHD VDDHD PCH L=60N W=600N M=1
MM5 N3 IN1A VDDHD VDDHD PCH L=60N W=600N M=1
MM25 N1 IN2 VDDHD VDDHD PCH L=60N W=600N M=2
MM24 N3 IN2 VDDHD VDDHD PCH L=60N W=600N M=2
MM23 N6 IN2 VDDHD VDDHD PCH L=60N W=600N M=2
MM22 N4 IN2 VDDHD VDDHD PCH L=60N W=600N M=2
MM18 N4 IN0A VDDHD VDDHD PCH L=60N W=600N M=1
MM17 N4 IN1B VDDHD VDDHD PCH L=60N W=600N M=1
MM16 N6 IN0B VDDHD VDDHD PCH L=60N W=600N M=1
MM15 N6 IN1B VDDHD VDDHD PCH L=60N W=600N M=1
XINV0 N1 VSSI VDDHD PREDEC0 S1AHSF400W40_AINV FN=2 WN=0.2U LN=0.06U FP=2 WP=0.4U LP=0.06U 
+ M=1
XINV1 N3 VSSI VDDHD PREDEC1 S1AHSF400W40_AINV FN=2 WN=0.2U LN=0.06U FP=2 WP=0.4U LP=0.06U 
+ M=1
XINV2 N4 VSSI VDDHD PREDEC2 S1AHSF400W40_AINV FN=2 WN=0.2U LN=0.06U FP=2 WP=0.4U LP=0.06U 
+ M=1
XINV3 N6 VSSI VDDHD PREDEC3 S1AHSF400W40_AINV FN=2 WN=0.2U LN=0.06U FP=2 WP=0.4U LP=0.06U 
+ M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CKBUF_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CKBUF_SB CK1B CK2 CKP CLK VDDHD VSSI
*.PININFO CKP:I CLK:I CK1B:O CK2:O VDDHD:B VSSI:B
XI28 CKP CLK VSSI VDDHD CK1B S1AHSF400W40_ANOR FN2=5 WN2=0.8U LN2=0.06U FN1=5 WN1=0.8U 
+ LN1=0.06U FP1=5 WP1=3U LP1=0.06U FP2=5 WP2=3U LP2=0.06U M=1
XINV0 CK1B VSSI VDDHD CK2 S1AHSF400W40_AINV FN=3 WN=0.7U LN=0.06U FP=3 WP=1.3U LP=0.06U 
+ M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    DECB1_X2_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_DECB1_X2_SB CLK CLK_ENV DEC EN ENC PD PREDEC VDDHD VSSI
*.PININFO CLK:I CLK_ENV:I EN:I ENC:I PD:I PREDEC:I DEC:O VDDHD:B VSSI:B
MM5 DEC PD VSSI VSSI NCH L=60N W=300N M=1
MM8 NT1 PREDEC ENC VSSI NCH L=60N W=1.5U M=2
MN0 DEC NT1 VSSI VSSI NCH L=60N W=1.25U M=4
MM6 NT1 EN VDDHD VDDHD PCH L=60N W=800N M=2
MM4 NT1 PREDEC VDDHD VDDHD PCH L=60N W=500N M=1
MM2 CLK_ENV CLK NT1 VDDHD PCH L=60N W=250.0N M=2
MP0 DEC NT1 VDDHD VDDHD PCH L=60N W=2.5U M=4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CDEC_M8_882_BIST_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CDEC_M8_882_BIST_SB BIST1B BIST2 BLEQ CEB CEBM CK1B CK2 CKD CKP CKPD 
+ CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN PD RE RSC VDDHD VDDI VSSI WE WEBXL 
+ WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] XM[0] XM[1] XM[2] XM[3] XM[4] 
+ XM[5] XM[6] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3] AX[0] 
+ AX[1] AX[2] AX[3] AX[4] AX[5] AX[6]
*.PININFO BIST1B:I BIST2:I CEB:I CEBM:I CKP:I CKPD:I CLK:I PD:I RSC:I WEBXL:I 
*.PININFO WEBXL1B:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I XM[0]:I 
*.PININFO XM[1]:I XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I Y[0]:I Y[1]:I Y[2]:I 
*.PININFO Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I BLEQ:O CK1B:O CK2:O CKD:O 
*.PININFO DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O 
*.PININFO DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O 
*.PININFO DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O 
*.PININFO DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O 
*.PININFO DEC_Y[3]:O DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O EN:O RE:O 
*.PININFO WE:O YL[0]:O YL[1]:O AX[0]:O AX[1]:O AX[2]:O AX[3]:O AX[4]:O AX[5]:O 
*.PININFO AX[6]:O VDDHD:B VDDI:B VSSI:B
XIPDEC_X0<0> AXC[0] AXT[0] AXC[1] AXT[1] AXC[2] PD DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] VDDHD VSSI S1AHSF400W40_DECB4_882_SB
XIPDEC_X0<1> AXC[0] AXT[0] AXC[1] AXT[1] AXT[2] PD DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] VDDHD VSSI S1AHSF400W40_DECB4_882_SB
XIPDEC_X1<0> AXC[3] AXT[3] AXC[4] AXT[4] AXC[5] PD DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] VDDHD VSSI S1AHSF400W40_DECB4_882_SB
XIPDEC_X1<1> AXC[3] AXT[3] AXC[4] AXT[4] AXT[5] PD DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] VDDHD VSSI S1AHSF400W40_DECB4_882_SB
XCEBBUF BIST1B BIST2 CEB CEBM CK1B CK2 CKPD CLK CLK_ENV EN ENC RSC VDDHD VSSI 
+ S1AHSF400W40_ENBUFB_BIST_SB
XABUF_Y<3> Y[3] YM[3] NET206 AYC[3] AYT[3] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<0> X[0] XM[0] AX[0] AXC[0] AXT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<1> X[1] XM[1] AX[1] AXC[1] AXT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<2> X[2] XM[2] AX[2] AXC[2] AXT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_Y<2> Y[2] YM[2] NET228 AYC[2] AYT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<6> X[6] XM[6] AX[6] AXC[6] AXT[6] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<3> X[3] XM[3] AX[3] AXC[3] AXT[3] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<4> X[4] XM[4] AX[4] AXC[4] AXT[4] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<5> X[5] XM[5] AX[5] AXC[5] AXT[5] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_Y<0> Y[0] YM[0] NET258[0] AYC[0] AYT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_Y<1> Y[1] YM[1] NET258[1] AYC[1] AYT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XIDEC_Y<4> NET024 NET024 DEC_Y[4] NET024 NET024 PD XY[4] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<5> NET024 NET024 DEC_Y[5] NET024 NET024 PD XY[5] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<6> NET024 NET024 DEC_Y[6] NET024 NET024 PD XY[6] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<7> NET024 NET024 DEC_Y[7] NET024 NET024 PD XY[7] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<0> NET0253 NET0253 DEC_Y[0] NET0253 NET0253 PD XY[0] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<1> NET0253 NET0253 DEC_Y[1] NET0253 NET0253 PD XY[1] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<2> NET0253 NET0253 DEC_Y[2] NET0253 NET0253 PD XY[2] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<3> NET0253 NET0253 DEC_Y[3] NET0253 NET0253 PD XY[3] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XDECB1_BLEQ BLEQ CKPD CLK_ENV ENC EN PD VDDHD VDDI VSSI S1AHSF400W40_DECB1_BLEQ_SB
XPREDEC_Y<0> AYC[0] AYT[0] AYC[1] AYT[1] AYC[2] XY[0] XY[1] XY[2] XY[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XPREDEC_Y<1> AYC[0] AYT[0] AYC[1] AYT[1] AYT[2] XY[4] XY[5] XY[6] XY[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XCKBUF CK1B CK2 CKP CLK VDDHD VSSI S1AHSF400W40_CKBUF_SB
XIDEC_CKD CLK CLK_ENV CKD EN ENC PD WEBXL1B VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_REWE<0> CLK CLK_ENV RE EN ENC PD WEBXL VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_REWE<1> CLK CLK_ENV WE EN ENC PD WEBXL1B VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_YL<0> CLK CLK_ENV YL[0] EN ENC PD AYC[3] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_YL<1> CLK CLK_ENV YL[1] EN ENC PD AYT[3] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<0> CLK CLK_ENV DEC_X2[0] EN ENC PD AXC[6] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<1> CLK CLK_ENV DEC_X2[1] EN ENC PD AXT[6] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_882_BIST_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_882_BIST_SB AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM 
+ CKD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE 
+ TK TM TRKBL VDDHD VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] 
+ X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] 
+ XM[5] XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] 
+ YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I RTSEL[0]:I RTSEL[1]:I 
*.PININFO TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I 
*.PININFO X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I XM[0]:I XM[1]:I 
*.PININFO XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I Y[0]:I 
*.PININFO Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O 
*.PININFO BIST2IO:O BLEQ:O BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O 
*.PININFO DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O 
*.PININFO DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O 
*.PININFO DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O DEC_X2[5]:O 
*.PININFO DEC_X2[6]:O DEC_X2[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O 
*.PININFO DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O PD_BUF:O RE:O SAE:O 
*.PININFO VHI:O VLO:O WE:O YL[0]:O YL[1]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B
XCOTHERS AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKP CKPD CLK 
+ DEC_X2[0] DEC_X2[1] EN PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL 
+ VDDHD VDDI VHI VLO VSSI WEB WEBM WEBXL WEBXL1B SAE WLP_SAEB NET95 WTSEL[0] 
+ WTSEL[1] WTSEL[2] S1AHSF400W40_COTH_BIST_882_SB
XCDEC BIST1B BIST2 BLEQ CEB CEBM CK1B CK2 CKD CKP CKPD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] EN PD_BUF RE RSC VDDHD VDDI VSSI WE WEBXL WEBXL1B X[0] 
+ X[1] X[2] X[3] X[4] X[5] X[6] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] Y[0] 
+ Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3] AX[0] AX[1] AX[2] AX[3] 
+ AX[4] AX[5] AX[6] S1AHSF400W40_CDEC_M8_882_BIST_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_882_BIST_M4_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_882_BIST_M4_SB AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM 
+ CKD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE 
+ TK TM TRKBL VDDHD VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] 
+ X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] 
+ XM[5] XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] 
+ YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I RTSEL[0]:I RTSEL[1]:I 
*.PININFO TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I 
*.PININFO X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I XM[0]:I XM[1]:I 
*.PININFO XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I Y[0]:I 
*.PININFO Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O 
*.PININFO BIST2IO:O BLEQ:O BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O 
*.PININFO DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O 
*.PININFO DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O 
*.PININFO DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O DEC_X2[5]:O 
*.PININFO DEC_X2[6]:O DEC_X2[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O 
*.PININFO DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O PD_BUF:O RE:O SAE:O 
*.PININFO VHI:O VLO:O WE:O YL[0]:O YL[1]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B
XCNT AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] 
+ DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] 
+ DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] 
+ DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] DEC_X2[5] 
+ DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] 
+ X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] 
+ XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3] 
+ S1AHSF400W40_CNT_CORE_882_BIST_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_882_BIST_M8M16_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_882_BIST_M8M16_SB AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB 
+ CEBM CKD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE 
+ TK TM TRKBL VDDHD VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] 
+ X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] 
+ XM[5] XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] 
+ YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I RTSEL[0]:I RTSEL[1]:I 
*.PININFO TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I 
*.PININFO X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I XM[0]:I XM[1]:I 
*.PININFO XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I Y[0]:I 
*.PININFO Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O 
*.PININFO BIST2IO:O BLEQ:O BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O 
*.PININFO DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O 
*.PININFO DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O 
*.PININFO DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O DEC_X2[5]:O 
*.PININFO DEC_X2[6]:O DEC_X2[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O 
*.PININFO DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O PD_BUF:O RE:O SAE:O 
*.PININFO VHI:O VLO:O WE:O YL[0]:O YL[1]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B
XCNT AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] 
+ DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] 
+ DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] 
+ DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] DEC_X2[5] 
+ DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] 
+ X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] 
+ XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3] 
+ S1AHSF400W40_CNT_CORE_882_BIST_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    WEBBUF_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_WEBBUF_SB BIST1B BIST2 CKC CKT VDDHD VSSI WEB WEBM WEBXL WEBXL1B
*.PININFO BIST1B:I BIST2:I CKC:I CKT:I WEB:I WEBM:I WEBXL:O WEBXL1B:O VDDHD:B 
*.PININFO VSSI:B
MM20 WEBXL CKC NET0115 VDDHD PCH L=60N W=300N M=1
MM21 NET0115 WEBXL1B VDDHD VDDHD PCH L=60N W=300N M=1
MM16 N5 CKT VDDHD VDDHD PCH L=60N W=1U M=2
MM6 WEBXL WEBX N5 VDDHD PCH L=60N W=1U M=2
MM10 WEBX WEB VDDHD VDDHD PCH L=60N W=600N M=1
MM0 WEBXL WEBX N7 VSSI NCH L=60N W=1U M=2
MM19 WEBXL CKT NET076 VSSI NCH L=60N W=200N M=1
MM18 NET076 WEBXL1B VSSI VSSI NCH L=60N W=200N M=1
MM12 WEBX WEB VSSI VSSI NCH L=60N W=300N M=1
MM17 N7 CKC VSSI VSSI NCH L=60N W=1U M=2
XI25 WEBXL VSSI VDDHD WEBXL1B S1AHSF400W40_AINV FN=2 WN=0.55U LN=0.06U FP=2 WP=1U 
+ LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    COTH_882_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_COTH_882_SB AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKP 
+ CKPD CLK DEC_X2[0] DEC_X2[1] EN PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM 
+ TRKBL VDDHD VDDI VHI VLO VSSI WEB WEBM WEBXL WEBXL1B WLP_SAE WLP_SAEB 
+ WLP_SAE_TK WTSEL[0] WTSEL[1] WTSEL[2]
*.PININFO AWT:I BIST:I CK1B:I CK2:I CLK:I DEC_X2[0]:I DEC_X2[1]:I EN:I PD:I 
*.PININFO PTSEL:I RTSEL[0]:I RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I 
*.PININFO WTSEL[1]:I WTSEL[2]:I AWT2:O BIST1B:O BIST2:O BIST2IO:O BLTRKWLDRV:O 
*.PININFO CKP:O CKPD:O PD_BUF:O RSC:O VHI:O VLO:O WEBXL:O WEBXL1B:O WLP_SAE:O 
*.PININFO WLP_SAEB:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE_TK:B
XWEBBUF_SB BIST1B BIST2 CK1B CK2 VDDHD VSSI WEB WEBM WEBXL WEBXL1B S1AHSF400W40_WEBBUF_SB
XVHILO_SB VDDHD VHI VLO VSSI S1AHSF400W40_VHILO_SB
XCKG CKP CLK EN RSC RSTCK TM VDDHD VSSI S1AHSF400W40_CKG_882_SB
XRESETD BLTRKWLDRV CK2 CKP CKPD CKPDCLK DEC_X2[0] DEC_X2[1] WLP_SAEB RSTCK TK 
+ TRKBL VDDHD VSSI WEBXL WLP_SAE WLP_SAE_TK PTSEL RTSEL[0] RTSEL[1] WTSEL[0] 
+ WTSEL[1] WTSEL[2] S1AHSF400W40_RESETD_882_SB
XPDBUF_SB PD PD_BUF VDDI VSSI S1AHSF400W40_PDBUF_SB
MP1 VDDHD PD VDDI VDDI PCH L=60N W=3U M=9
MP0 VDDHD PD VDDI VDDI PCH L=60N W=3.8U M=16
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    ABUF_882_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ABUF_882_SB A AM AX1B AX1BL AX1BL1B BIST1B BIST2 CK1B CK2 VDDHD VSSI
*.PININFO A:I AM:I BIST1B:I BIST2:I CK1B:I CK2:I AX1B:O AX1BL:O AX1BL1B:O 
*.PININFO VDDHD:B VSSI:B
MM26 AX1BL CK1B NET57 VDDHD PCH L=60N W=300N M=1
MM28 N5 CK2 VDDHD VDDHD PCH L=60N W=1U M=4
MM27 NET57 AX1BL1B VDDHD VDDHD PCH L=60N W=300N M=1
MM29 AX1BL A N5 VDDHD PCH L=60N W=1U M=2
MM20 AX1BL CK2 NET82 VSSI NCH L=60N W=200N M=1
MM23 N7 CK1B VSSI VSSI NCH L=60N W=1U M=4
MM19 AX1BL A N7 VSSI NCH L=60N W=1U M=2
MM21 NET82 AX1BL1B VSSI VSSI NCH L=60N W=200N M=1
XI25 AX1BL VSSI VDDHD AX1BL1B S1AHSF400W40_AINV FN=2 WN=0.55U LN=0.06U FP=2 WP=1U 
+ LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    ABUF_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ABUF_SB A AM AX1B AX1BL AX1BL1B BIST1B BIST2 CK1B CK2 VDDHD VSSI
*.PININFO A:I AM:I BIST1B:I BIST2:I CK1B:I CK2:I AX1B:O AX1BL:O AX1BL1B:O 
*.PININFO VDDHD:B VSSI:B
MM26 AX1BL CK1B NET57 VDDHD PCH L=60N W=300N M=1
MM28 N5 CK2 VDDHD VDDHD PCH L=60N W=1U M=2
MM27 NET57 AX1BL1B VDDHD VDDHD PCH L=60N W=300N M=1
MM29 AX1BL A N5 VDDHD PCH L=60N W=1U M=2
MM20 AX1BL CK2 NET82 VSSI NCH L=60N W=200N M=1
MM23 N7 CK1B VSSI VSSI NCH L=60N W=1U M=2
MM19 AX1BL A N7 VSSI NCH L=60N W=1U M=2
MM21 NET82 AX1BL1B VSSI VSSI NCH L=60N W=200N M=1
XI25 AX1BL VSSI VDDHD AX1BL1B S1AHSF400W40_AINV FN=1 WN=0.55U LN=0.06U FP=1 WP=1U 
+ LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    ENBUFB_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ENBUFB_SB BIST1B BIST2 CEB CEBM CK1B CK2 CKP CLK CLK_ENV EN ENC RSC 
+ VDDHD VSSI
*.PININFO BIST1B:I BIST2:I CEB:I CEBM:I CK1B:I CK2:I CKP:I CLK:I RSC:I 
*.PININFO CLK_ENV:O EN:O ENC:O VDDHD:B VSSI:B
XI141 CEBXL VSSI VDDHD EN S1AHSF400W40_AINV FN=3 WN=1U LN=0.06U FP=3 WP=2U LP=0.06U M=1
MM18 N7 CK1B NET120 VSSI NCH L=60N W=1U M=1
MM17 CEBXL CEBX N7 VSSI NCH L=60N W=1U M=1
MM3 CEBXL CK2 NET112 VSSI NCH L=60N W=500N M=1
MM4 NET112 EN NET108 VSSI NCH L=60N W=500N M=1
MM20 NET120 RSC VSSI VSSI NCH L=60N W=1U M=2
MM22 ENC CLK NET143 VSSI NCH L=60N W=3.2U M=5
MM12 CEBX CEB VSSI VSSI NCH L=60N W=500N M=1
MM5 NET108 RSC VSSI VSSI NCH L=60N W=1U M=1
MM23 ENC CKP NET143 VSSI NCH L=60N W=3.2U M=1
MM0 NET143 EN VSSI VSSI NCH L=60N W=3.2U M=5
MM1 CEBXL CK1B NET179 VDDHD PCH L=60N W=500N M=1
MM10 CEBX CEB VDDHD VDDHD PCH L=60N W=500N M=1
MM19 N5 CK2 VDDHD VDDHD PCH L=60N W=1U M=2
MM16 CEBXL CEBX N5 VDDHD PCH L=60N W=1U M=2
MM7 CEBXL RSC VDDHD VDDHD PCH L=60N W=700N M=2
MM21 VDDHD EN ENC VDDHD PCH L=60N W=700N M=3
MM6 VDDHD CKP CLK_ENV VDDHD PCH L=60N W=750.0N M=4
MM2 NET179 EN VDDHD VDDHD PCH L=60N W=500N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CDEC_M8_882_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CDEC_M8_882_SB BIST1B BIST2 BLEQ CEB CEBM CK1B CK2 CKD CKP CKPD CLK 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN PD RE RSC VDDHD VDDI VSSI WE WEBXL 
+ WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] XM[0] XM[1] XM[2] XM[3] XM[4] 
+ XM[5] XM[6] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3] AX[0] 
+ AX[1] AX[2] AX[3] AX[4] AX[5] AX[6]
*.PININFO BIST1B:I BIST2:I CEB:I CEBM:I CKP:I CKPD:I CLK:I PD:I RSC:I WEBXL:I 
*.PININFO WEBXL1B:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I XM[0]:I 
*.PININFO XM[1]:I XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I Y[0]:I Y[1]:I Y[2]:I 
*.PININFO Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I BLEQ:O CK1B:O CK2:O CKD:O 
*.PININFO DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O 
*.PININFO DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O 
*.PININFO DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O 
*.PININFO DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O 
*.PININFO DEC_Y[3]:O DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O EN:O RE:O 
*.PININFO WE:O YL[0]:O YL[1]:O AX[0]:O AX[1]:O AX[2]:O AX[3]:O AX[4]:O AX[5]:O 
*.PININFO AX[6]:O VDDHD:B VDDI:B VSSI:B
XABUF_X<6> X[6] XM[6] AX[6] AXC[6] AXT[6] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_882_SB
XIPDEC_X0<0> AXC[0] AXT[0] AXC[1] AXT[1] AXC[2] PD DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] VDDHD VSSI S1AHSF400W40_DECB4_882_SB
XIPDEC_X0<1> AXC[0] AXT[0] AXC[1] AXT[1] AXT[2] PD DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] VDDHD VSSI S1AHSF400W40_DECB4_882_SB
XIPDEC_X1<0> AXC[3] AXT[3] AXC[4] AXT[4] AXC[5] PD DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] VDDHD VSSI S1AHSF400W40_DECB4_882_SB
XIPDEC_X1<1> AXC[3] AXT[3] AXC[4] AXT[4] AXT[5] PD DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] VDDHD VSSI S1AHSF400W40_DECB4_882_SB
XIDEC_Y<4> NET024 NET024 DEC_Y[4] NET024 NET024 PD XY[4] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<5> NET024 NET024 DEC_Y[5] NET024 NET024 PD XY[5] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<6> NET024 NET024 DEC_Y[6] NET024 NET024 PD XY[6] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<7> NET024 NET024 DEC_Y[7] NET024 NET024 PD XY[7] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<0> NET0253 NET0253 DEC_Y[0] NET0253 NET0253 PD XY[0] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<1> NET0253 NET0253 DEC_Y[1] NET0253 NET0253 PD XY[1] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<2> NET0253 NET0253 DEC_Y[2] NET0253 NET0253 PD XY[2] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<3> NET0253 NET0253 DEC_Y[3] NET0253 NET0253 PD XY[3] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XDECB1_BLEQ BLEQ CKPD CLK_ENV ENC EN PD VDDHD VDDI VSSI S1AHSF400W40_DECB1_BLEQ_SB
XPREDEC_Y<0> AYC[0] AYT[0] AYC[1] AYT[1] AYC[2] XY[0] XY[1] XY[2] XY[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XPREDEC_Y<1> AYC[0] AYT[0] AYC[1] AYT[1] AYT[2] XY[4] XY[5] XY[6] XY[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XCKBUF CK1B CK2 CKP CLK VDDHD VSSI S1AHSF400W40_CKBUF_SB
XABUF_Y<3> Y[3] YM[3] NET206 AYC[3] AYT[3] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<0> X[0] XM[0] AX[0] AXC[0] AXT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<1> X[1] XM[1] AX[1] AXC[1] AXT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<2> X[2] XM[2] AX[2] AXC[2] AXT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_Y<2> Y[2] YM[2] NET228 AYC[2] AYT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<3> X[3] XM[3] AX[3] AXC[3] AXT[3] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<4> X[4] XM[4] AX[4] AXC[4] AXT[4] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<5> X[5] XM[5] AX[5] AXC[5] AXT[5] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_Y<0> Y[0] YM[0] NET258[0] AYC[0] AYT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_Y<1> Y[1] YM[1] NET258[1] AYC[1] AYT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XCEBBUF BIST1B BIST2 CEB CEBM CK1B CK2 CKPD CLK CLK_ENV EN ENC RSC VDDHD VSSI 
+ S1AHSF400W40_ENBUFB_SB
XIDEC_CKD CLK CLK_ENV CKD EN ENC PD WEBXL1B VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_REWE<0> CLK CLK_ENV RE EN ENC PD WEBXL VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_REWE<1> CLK CLK_ENV WE EN ENC PD WEBXL1B VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_YL<0> CLK CLK_ENV YL[0] EN ENC PD AYC[3] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_YL<1> CLK CLK_ENV YL[1] EN ENC PD AYT[3] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<0> CLK CLK_ENV DEC_X2[0] EN ENC PD AXC[6] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<1> CLK CLK_ENV DEC_X2[1] EN ENC PD AXT[6] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_882_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_882_SB AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM CKD CLK 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] 
+ DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE TK TM 
+ TRKBL VDDHD VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] X[0] 
+ X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I RTSEL[0]:I RTSEL[1]:I 
*.PININFO TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I 
*.PININFO X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I XM[0]:I XM[1]:I 
*.PININFO XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I Y[0]:I 
*.PININFO Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O 
*.PININFO BIST2IO:O BLEQ:O BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O 
*.PININFO DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O 
*.PININFO DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O 
*.PININFO DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O DEC_X2[5]:O 
*.PININFO DEC_X2[6]:O DEC_X2[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O 
*.PININFO DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O PD_BUF:O RE:O SAE:O 
*.PININFO VHI:O VLO:O WE:O YL[0]:O YL[1]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B
XCOTHERS AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKP CKPD CLK 
+ DEC_X2[0] DEC_X2[1] EN PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL 
+ VDDHD VDDI VHI VLO VSSI WEB WEBM WEBXL WEBXL1B SAE WLP_SAEB NET95 WTSEL[0] 
+ WTSEL[1] WTSEL[2] S1AHSF400W40_COTH_882_SB
XCDEC BIST1B BIST2 BLEQ CEB CEBM CK1B CK2 CKD CKP CKPD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] EN PD_BUF RE RSC VDDHD VDDI VSSI WE WEBXL WEBXL1B X[0] 
+ X[1] X[2] X[3] X[4] X[5] X[6] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] Y[0] 
+ Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3] AX[0] AX[1] AX[2] AX[3] 
+ AX[4] AX[5] AX[6] S1AHSF400W40_CDEC_M8_882_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_882_M4_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_882_M4_SB AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM CKD 
+ CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] 
+ DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE TK TM 
+ TRKBL VDDHD VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] X[0] 
+ X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I RTSEL[0]:I RTSEL[1]:I 
*.PININFO TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I 
*.PININFO X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I XM[0]:I XM[1]:I 
*.PININFO XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I Y[0]:I 
*.PININFO Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O 
*.PININFO BIST2IO:O BLEQ:O BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O 
*.PININFO DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O 
*.PININFO DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O 
*.PININFO DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O DEC_X2[5]:O 
*.PININFO DEC_X2[6]:O DEC_X2[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O 
*.PININFO DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O PD_BUF:O RE:O SAE:O 
*.PININFO VHI:O VLO:O WE:O YL[0]:O YL[1]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B
XCNT AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] 
+ DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] 
+ DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] 
+ DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] DEC_X2[5] 
+ DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] 
+ X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] 
+ XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3] 
+ S1AHSF400W40_CNT_CORE_882_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_882_M8M16_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_882_M8M16_SB AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM 
+ CKD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE 
+ TK TM TRKBL VDDHD VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] 
+ X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] 
+ XM[5] XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] 
+ YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I RTSEL[0]:I RTSEL[1]:I 
*.PININFO TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I 
*.PININFO X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I XM[0]:I XM[1]:I 
*.PININFO XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I Y[0]:I 
*.PININFO Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O 
*.PININFO BIST2IO:O BLEQ:O BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O 
*.PININFO DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O 
*.PININFO DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O 
*.PININFO DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O DEC_X2[5]:O 
*.PININFO DEC_X2[6]:O DEC_X2[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O 
*.PININFO DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O PD_BUF:O RE:O SAE:O 
*.PININFO VHI:O VLO:O WE:O YL[0]:O YL[1]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B
XCNT AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] 
+ DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] 
+ DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] 
+ DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] DEC_X2[5] 
+ DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] 
+ X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] 
+ XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3] 
+ S1AHSF400W40_CNT_CORE_882_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CKG_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CKG_SB CKP CLK EN RSC RSTCK TM VDDHD VSSI
*.PININFO CLK:I EN:I RSTCK:I TM:I CKP:O RSC:O VDDHD:B VSSI:B
XINV0 Z17 VSSI VDDHD RSC S1AHSF400W40_AINV FN=3 WN=0.35U LN=0.06U FP=3 WP=0.7U LP=0.06U 
+ M=1
XI50 RSTCK CKP VSSI VDDHD RSCI S1AHSF400W40_ANAND FN2=1 WN2=2U LN2=0.06U FN1=1 WN1=2U 
+ LN1=0.06U FP1=1 WP1=2U LP1=0.06U FP2=1 WP2=2U LP2=0.06U M=1
XNAND4 CKPC Z19 VSSI VDDHD CKP S1AHSF400W40_ANAND FN2=4 WN2=0.75U LN2=0.06U FN1=4 
+ WN1=0.75U LN1=0.06U FP1=4 WP1=3U LP1=0.06U FP2=4 WP2=1.5U LP2=0.06U M=1
XNAND5 CKP RSC VSSI VDDHD Z19 S1AHSF400W40_ANAND FN2=1 WN2=0.54U LN2=0.06U FN1=1 
+ WN1=0.54U LN1=0.06U FP1=1 WP1=0.75U LP1=0.06U FP2=1 WP2=0.75U LP2=0.06U M=1
XNAND3 Z16 Z14 VSSI VDDHD Z17 S1AHSF400W40_ANAND FN2=1 WN2=0.54U LN2=0.06U FN1=1 
+ WN1=0.54U LN1=0.06U FP1=1 WP1=0.54U LP1=0.06U FP2=1 WP2=0.54U LP2=0.06U M=1
XI49 Z17 CLK VSSI VDDHD Z14 S1AHSF400W40_ANAND FN2=1 WN2=0.4U LN2=0.06U FN1=1 WN1=0.4U 
+ LN1=0.06U FP1=1 WP1=0.4U LP1=0.06U FP2=1 WP2=0.4U LP2=0.06U M=1
XNAND0 TM CLK VSSI VDDHD Z15 S1AHSF400W40_ANAND FN2=1 WN2=0.4U LN2=0.06U FN1=1 WN1=0.4U 
+ LN1=0.06U FP1=1 WP1=0.4U LP1=0.06U FP2=1 WP2=0.4U LP2=0.06U M=1
XNAND12 CLK RSC EN VSSI VDDHD CKPC S1AHSF400W40_ANAND3 FN3=1 WN3=2U LN3=0.06U FN2=1 
+ WN2=2U LN2=0.06U FN1=1 WN1=2U LN1=0.06U FP1=1 WP1=1U LP1=0.06U FP2=1 WP2=1U 
+ LP2=0.06U FP3=1 WP3=1U LP3=0.06U M=1
XI53 RSTCK CKP Z15 VSSI VDDHD Z16 S1AHSF400W40_ANAND3 FN3=1 WN3=0.9U LN3=0.06U FN2=1 
+ WN2=0.9U LN2=0.06U FN1=1 WN1=0.9U LN1=0.06U FP1=1 WP1=0.6U LP1=0.06U FP2=1 
+ WP2=0.6U LP2=0.06U FP3=1 WP3=0.6U LP3=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    RESETD_WTSEL_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_RESETD_WTSEL_SB CKP V[0] V[1] VDDHD VSSI TD_01_11 TD_10
*.PININFO CKP:I V[0]:I V[1]:I TD_01_11:O TD_10:O VDDHD:B VSSI:B
XI21 CKP VSSI VDDHD Z0 S1AHSF400W40_AINV FN=1 WN=0.3U LN=180N FP=1 WP=0.6U LP=180N M=1
XI76 Z0 V[0] VSSI VDDHD TD_01_11 S1AHSF400W40_ANAND FN2=1 WN2=0.6U LN2=0.18U FN1=1 
+ WN1=0.6U LN1=0.18U FP1=1 WP1=0.6U LP1=0.18U FP2=1 WP2=0.6U LP2=0.18U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    RESETD_RTSEL_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_RESETD_RTSEL_SB CKP V[0] V[1] VDDHD VSSI TD_01_11 TD_10
*.PININFO CKP:I V[0]:I V[1]:I TD_01_11:O TD_10:O VDDHD:B VSSI:B
XI21 CKP VSSI VDDHD Z3 S1AHSF400W40_AINV FN=1 WN=0.3U LN=180N FP=1 WP=0.6U LP=180N M=1
XI78 Z4 VSSI VDDHD Z5 S1AHSF400W40_AINV FN=1 WN=0.3U LN=180N FP=1 WP=0.6U LP=180N M=1
XI77 Z3 VSSI VDDHD Z4 S1AHSF400W40_AINV FN=1 WN=0.3U LN=180N FP=1 WP=0.6U LP=180N M=1
XND0 CKP TD_10 VSSI VDDHD Z0 S1AHSF400W40_ANAND FN2=1 WN2=0.6U LN2=0.06U FN1=1 WN1=0.6U 
+ LN1=0.06U FP1=1 WP1=0.6U LP1=0.06U FP2=1 WP2=0.6U LP2=0.06U M=1
XI76 Z0 V[0] VSSI VDDHD TD_01_11 S1AHSF400W40_ANAND FN2=1 WN2=0.6U LN2=0.06U FN1=1 
+ WN1=0.6U LN1=0.06U FP1=1 WP1=0.6U LP1=0.06U FP2=1 WP2=0.6U LP2=0.06U M=1
XI79 Z5 V[1] VSSI VDDHD TD_10 S1AHSF400W40_ANAND FN2=1 WN2=0.6U LN2=0.18U FN1=1 WN1=0.6U 
+ LN1=0.18U FP1=1 WP1=0.6U LP1=0.18U FP2=1 WP2=0.6U LP2=0.18U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    RESETD_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_RESETD_SB BLTRKWLDRV CK2 CKP CKPD CKPDCLK IOSAEB RSTCK TK TRKBL VDDHD 
+ VSSI WEBXL WLP_SAE WLP_SAE_TK PTSEL RV[0] RV[1] WV[0] WV[1] WV[2]
*.PININFO CK2:I CKP:I WEBXL:I PTSEL:I RV[0]:I RV[1]:I WV[0]:I WV[1]:I WV[2]:I 
*.PININFO BLTRKWLDRV:O CKPD:O CKPDCLK:O IOSAEB:O RSTCK:O WLP_SAE:O TK:B 
*.PININFO TRKBL:B VDDHD:B VSSI:B WLP_SAE_TK:B
XTSEL_WT TRKBL1B WV[0] WV[1] VDDHD VSSI NET118 NET115 S1AHSF400W40_RESETD_WTSEL_SB
XTSEL_RT CKP RV[0] RV[1] VDDHD VSSI RTD_01_11 RTD_10 S1AHSF400W40_RESETD_RTSEL_SB
XI668 SHORT_D1 VSSI VDDHD NET0145 S1AHSF400W40_AINV FN=1 WN=0.4U LN=60N FP=1 WP=0.8U 
+ LP=60N M=1
XI653 SAE_FIRE2 VSSI VDDHD WLP_SAE S1AHSF400W40_AINV FN=12 WN=0.5U LN=60N FP=6 WP=2U 
+ LP=60N M=1
XI537 RTKB2 VSSI VDDHD BLTRKWLDRV S1AHSF400W40_AINV FN=12 WN=0.5U LN=60N FP=6 WP=2U 
+ LP=60N M=1
XI593 CKP VSSI VDDHD Z1 S1AHSF400W40_AINV FN=1 WN=1U LN=0.06U FP=1 WP=2U LP=0.06U M=1
XI594 Z1 VSSI VDDHD CKPD S1AHSF400W40_AINV FN=8 WN=0.5U LN=0.06U FP=4 WP=2U LP=0.06U M=1
XI661 TRKBL1B VSSI VDDHD TRKBL2 S1AHSF400W40_AINV FN=2 WN=0.25U LN=60N FP=2 WP=0.5U 
+ LP=60N M=1
XI540 RTKB1B VSSI VDDHD RTKB2 S1AHSF400W40_AINV FN=6 WN=0.4U LN=60N FP=6 WP=0.8U LP=60N 
+ M=1
XI541 RTKB VSSI VDDHD RTKB1B S1AHSF400W40_AINV FN=2 WN=0.4U LN=60N FP=2 WP=0.8U LP=60N M=1
XI574 TRKBL VSSI VDDHD TRKBL1B S1AHSF400W40_AINV FN=3 WN=0.35U LN=90N FP=3 WP=0.7U LP=90N 
+ M=1
XI669 NET0145 VSSI VDDHD SHORT_D2 S1AHSF400W40_AINV FN=1 WN=0.4U LN=60N FP=1 WP=0.8U 
+ LP=60N M=1
XI675 TRKBL1B NET118 VSSI VDDHD NET0187 S1AHSF400W40_ANAND FN2=1 WN2=0.6U LN2=60N FN1=1 
+ WN1=0.6U LN1=60N FP1=1 WP1=0.6U LP1=60N FP2=1 WP2=0.6U LP2=60N M=1
XI666 SHORT_D2 TRKBL2 VSSI VDDHD TRKBL2B S1AHSF400W40_ANAND FN2=2 WN2=0.5U LN2=90N FN1=2 
+ WN1=0.5U LN1=60N FP1=2 WP1=0.5U LP1=60N FP2=2 WP2=0.5U LP2=90N M=1
XI658 WV[2] RTKB1B VSSI VDDHD SHORT_D1 S1AHSF400W40_ANAND FN2=1 WN2=0.6U LN2=60N FN1=1 
+ WN1=0.6U LN1=60N FP1=1 WP1=0.6U LP1=60N FP2=1 WP2=0.6U LP2=60N M=1
XI654 SHORT_D1 NET0187 VSSI VDDHD RSTCK S1AHSF400W40_ANAND FN2=2 WN2=0.75U LN2=60N FN1=2 
+ WN1=0.75U LN1=60N FP1=2 WP1=0.75U LP1=60N FP2=2 WP2=0.75U LP2=60N M=1
XI667 WEBXL BLTRKWLDRV TRKBL2B VSSI VDDHD SAE_FIRE2 S1AHSF400W40_ANAND3 FN3=1 WN3=3U 
+ LN3=60N FN2=1 WN2=3U LN2=60N FN1=1 WN1=3U LN1=60N FP1=1 WP1=3U LP1=60N FP2=1 
+ WP2=3U LP2=60N FP3=1 WP3=3U LP3=60N M=1
XI584 CKP RTD_01_11 RTD_10 VSSI VDDHD RTKB S1AHSF400W40_ANAND3 FN3=2 WN3=0.6U LN3=60N 
+ FN2=2 WN2=0.6U LN2=60N FN1=2 WN1=0.6U LN1=60N FP1=2 WP1=0.4U LP1=60N FP2=2 
+ WP2=0.4U LP2=60N FP3=2 WP3=0.4U LP3=60N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    COTH_BIST_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_COTH_BIST_SB AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 
+ CKP CKPD CLK EN PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL VDDHD VDDI 
+ VHI VLO VSSI WEB WEBM WEBXL WEBXL1B WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] 
+ WTSEL[1] WTSEL[2]
*.PININFO AWT:I BIST:I CK1B:I CK2:I CLK:I EN:I PD:I PTSEL:I RTSEL[0]:I 
*.PININFO RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I AWT2:O 
*.PININFO BIST1B:O BIST2:O BIST2IO:O BLTRKWLDRV:O CKP:O CKPD:O PD_BUF:O RSC:O 
*.PININFO VHI:O VLO:O WEBXL:O WEBXL1B:O WLP_SAE:O WLP_SAEB:O TK:B TRKBL:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE_TK:B
MP1 VDDHD PD VDDI VDDI PCH L=60N W=3U M=22
MP0 VDDHD PD VDDI VDDI PCH L=60N W=3.8U M=29
XWEBBUF BIST1B BIST2 CK1B CK2 VDDHD VSSI WEB WEBM WEBXL WEBXL1B 
+ S1AHSF400W40_WEBBUF_BIST_SB
XVHILO_SB VDDHD VHI VLO VSSI S1AHSF400W40_VHILO_SB
XBISTD_SB BIST BIST1B BIST2 BIST2IO VDDHD VSSI S1AHSF400W40_BISTD_SB
XPDBUF_SB PD PD_BUF VDDI VSSI S1AHSF400W40_PDBUF_SB
XCKG CKP CLK EN RSC RSTCK TM VDDHD VSSI S1AHSF400W40_CKG_SB
XRESETD BLTRKWLDRV CK2 CKP CKPD CKPDCLK WLP_SAEB RSTCK TK TRKBL VDDHD VSSI 
+ WEBXL WLP_SAE WLP_SAE_TK PTSEL RTSEL[0] RTSEL[1] WTSEL[0] WTSEL[1] WTSEL[2] 
+ S1AHSF400W40_RESETD_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    DECB2_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_DECB2_SB IN0A IN0B IN1 PREDEC0 PREDEC1 VDDHD VSSI
*.PININFO IN0A:I IN0B:I IN1:I PREDEC0:O PREDEC1:O VDDHD:B VSSI:B
MM5 N3 IN1 VDDHD VDDHD PCH L=60N W=600N M=2
MM2 N1 IN1 VDDHD VDDHD PCH L=60N W=600N M=2
MM1 N1 IN0A VDDHD VDDHD PCH L=60N W=600N M=1
MM4 N3 IN0B VDDHD VDDHD PCH L=60N W=600N M=1
MM8 N2 IN1 VSSI VSSI NCH L=60N W=600N M=2
MM7 N3 IN0B N2 VSSI NCH L=60N W=600N M=1
MM0 N1 IN0A N2 VSSI NCH L=60N W=600N M=1
XINV0 N3 VSSI VDDHD PREDEC1 S1AHSF400W40_AINV FN=2 WN=0.2U LN=0.06U FP=2 WP=0.4U LP=0.06U 
+ M=1
XINV1 N1 VSSI VDDHD PREDEC0 S1AHSF400W40_AINV FN=2 WN=0.2U LN=0.06U FP=2 WP=0.4U LP=0.06U 
+ M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CDEC_M8_884_BIST_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CDEC_M8_884_BIST_SB BIST1B BIST2 BLEQ CEB CEBM CK1B CK2 CKD CKP CKPD 
+ CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_Y[0] 
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN PD RE RSC 
+ VDDHD VDDI VSSI WE WEBXL WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] 
+ XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] Y[0] Y[1] Y[2] Y[3] YL[0] 
+ YL[1] YM[0] YM[1] YM[2] YM[3] AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7]
*.PININFO BIST1B:I BIST2:I CEB:I CEBM:I CKP:I CKPD:I CLK:I PD:I RSC:I WEBXL:I 
*.PININFO WEBXL1B:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I 
*.PININFO Y[0]:I Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I BLEQ:O 
*.PININFO CK1B:O CK2:O CKD:O DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O 
*.PININFO DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O DEC_X1[0]:O 
*.PININFO DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O DEC_X1[5]:O 
*.PININFO DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O DEC_X2[2]:O 
*.PININFO DEC_X2[3]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O 
*.PININFO DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O EN:O RE:O WE:O YL[0]:O YL[1]:O 
*.PININFO AX[0]:O AX[1]:O AX[2]:O AX[3]:O AX[4]:O AX[5]:O AX[6]:O AX[7]:O 
*.PININFO VDDHD:B VDDI:B VSSI:B
XCEBBUF BIST1B BIST2 CEB CEBM CK1B CK2 CKPD CLK CLK_ENV EN ENC RSC VDDHD VSSI 
+ S1AHSF400W40_ENBUFB_BIST_SB
XABUF_Y<3> Y[3] YM[3] NET206 AYC[3] AYT[3] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<0> X[0] XM[0] AX[0] AXC[0] AXT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<1> X[1] XM[1] AX[1] AXC[1] AXT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<2> X[2] XM[2] AX[2] AXC[2] AXT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_Y<2> Y[2] YM[2] NET228 AYC[2] AYT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<6> X[6] XM[6] AX[6] AXC[6] AXT[6] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<7> X[7] XM[7] AX[7] AXC[7] AXT[7] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<3> X[3] XM[3] AX[3] AXC[3] AXT[3] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<4> X[4] XM[4] AX[4] AXC[4] AXT[4] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<5> X[5] XM[5] AX[5] AXC[5] AXT[5] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_Y<0> Y[0] YM[0] NET258[0] AYC[0] AYT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_Y<1> Y[1] YM[1] NET258[1] AYC[1] AYT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XIPDEC_X2<0> AXC[6] AXT[6] AXC[7] XC[0] XC[1] VDDHD VSSI S1AHSF400W40_DECB2_SB
XIPDEC_X2<1> AXC[6] AXT[6] AXT[7] XC[2] XC[3] VDDHD VSSI S1AHSF400W40_DECB2_SB
XIDEC_Y<0> NET0260 NET0260 DEC_Y[0] NET0260 NET0260 PD XY[0] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<1> NET0260 NET0260 DEC_Y[1] NET0260 NET0260 PD XY[1] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<2> NET0260 NET0260 DEC_Y[2] NET0260 NET0260 PD XY[2] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<3> NET0260 NET0260 DEC_Y[3] NET0260 NET0260 PD XY[3] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<4> NET0261 NET0261 DEC_Y[4] NET0261 NET0261 PD XY[4] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<5> NET0261 NET0261 DEC_Y[5] NET0261 NET0261 PD XY[5] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<6> NET0261 NET0261 DEC_Y[6] NET0261 NET0261 PD XY[6] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<7> NET0261 NET0261 DEC_Y[7] NET0261 NET0261 PD XY[7] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<0> NET0252 NET0252 DEC_X1[0] NET0252 NET0252 PD XB[0] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<1> NET0252 NET0252 DEC_X1[1] NET0252 NET0252 PD XB[1] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<2> NET0252 NET0252 DEC_X1[2] NET0252 NET0252 PD XB[2] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<3> NET0252 NET0252 DEC_X1[3] NET0252 NET0252 PD XB[3] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<4> NET0252 NET0252 DEC_X1[4] NET0252 NET0252 PD XB[4] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<5> NET0252 NET0252 DEC_X1[5] NET0252 NET0252 PD XB[5] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<6> NET0252 NET0252 DEC_X1[6] NET0252 NET0252 PD XB[6] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<7> NET0252 NET0252 DEC_X1[7] NET0252 NET0252 PD XB[7] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<0> NET0251 NET0251 DEC_X0[0] NET0251 NET0251 PD XA[0] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<1> NET0251 NET0251 DEC_X0[1] NET0251 NET0251 PD XA[1] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<2> NET0251 NET0251 DEC_X0[2] NET0251 NET0251 PD XA[2] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<3> NET0251 NET0251 DEC_X0[3] NET0251 NET0251 PD XA[3] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<4> NET0251 NET0251 DEC_X0[4] NET0251 NET0251 PD XA[4] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<5> NET0251 NET0251 DEC_X0[5] NET0251 NET0251 PD XA[5] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<6> NET0251 NET0251 DEC_X0[6] NET0251 NET0251 PD XA[6] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<7> NET0251 NET0251 DEC_X0[7] NET0251 NET0251 PD XA[7] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XDECB1_BLEQ BLEQ CKPD CLK_ENV ENC EN PD VDDHD VDDI VSSI S1AHSF400W40_DECB1_BLEQ_SB
XIPDEC_X0<0> AXC[0] AXT[0] AXC[1] AXT[1] AXC[2] XA[0] XA[1] XA[2] XA[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XIPDEC_X0<1> AXC[0] AXT[0] AXC[1] AXT[1] AXT[2] XA[4] XA[5] XA[6] XA[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XIPDEC_X1<0> AXC[3] AXT[3] AXC[4] AXT[4] AXC[5] XB[0] XB[1] XB[2] XB[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XIPDEC_X1<1> AXC[3] AXT[3] AXC[4] AXT[4] AXT[5] XB[4] XB[5] XB[6] XB[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XPREDEC_Y<0> AYC[0] AYT[0] AYC[1] AYT[1] AYC[2] XY[0] XY[1] XY[2] XY[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XPREDEC_Y<1> AYC[0] AYT[0] AYC[1] AYT[1] AYT[2] XY[4] XY[5] XY[6] XY[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XCKBUF CK1B CK2 CKPD CLK VDDHD VSSI S1AHSF400W40_CKBUF_SB
XIDEC_CKD CLK CLK_ENV CKD EN ENC PD WEBXL1B VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_REWE<0> CLK CLK_ENV RE EN ENC PD WEBXL VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_REWE<1> CLK CLK_ENV WE EN ENC PD WEBXL1B VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_YL<0> CLK CLK_ENV YL[0] EN ENC PD AYC[3] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_YL<1> CLK CLK_ENV YL[1] EN ENC PD AYT[3] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<0> CLK CLK_ENV DEC_X2[0] EN ENC PD XC[0] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<1> CLK CLK_ENV DEC_X2[1] EN ENC PD XC[1] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<2> CLK CLK_ENV DEC_X2[2] EN ENC PD XC[2] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<3> CLK CLK_ENV DEC_X2[3] EN ENC PD XC[3] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_884_BIST_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_884_BIST_SB AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM 
+ CKD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE 
+ TK TM TRKBL VDDHD VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] 
+ X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] 
+ XM[5] XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] 
+ YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I RTSEL[0]:I RTSEL[1]:I 
*.PININFO TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I 
*.PININFO X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I XM[0]:I XM[1]:I 
*.PININFO XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I Y[0]:I 
*.PININFO Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O 
*.PININFO BIST2IO:O BLEQ:O BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O 
*.PININFO DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O 
*.PININFO DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O 
*.PININFO DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O DEC_X2[5]:O 
*.PININFO DEC_X2[6]:O DEC_X2[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O 
*.PININFO DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O PD_BUF:O RE:O SAE:O 
*.PININFO VHI:O VLO:O WE:O YL[0]:O YL[1]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B
XCOTHERS AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKP CKPD CLK 
+ EN PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL VDDHD VDDI VHI VLO VSSI 
+ WEB WEBM WEBXL WEBXL1B SAE WLP_SAEB NET95 WTSEL[0] WTSEL[1] WTSEL[2] 
+ S1AHSF400W40_COTH_BIST_SB
XCDEC BIST1B BIST2 BLEQ CEB CEBM CK1B CK2 CKD CKP CKPD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN PD_BUF RE RSC VDDHD VDDI VSSI WE 
+ WEBXL WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] XM[0] XM[1] XM[2] 
+ XM[3] XM[4] XM[5] XM[6] XM[7] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] 
+ YM[2] YM[3] AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] 
+ S1AHSF400W40_CDEC_M8_884_BIST_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_884_BIST_M4_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_884_BIST_M4_SB AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM 
+ CKD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE 
+ TK TM TRKBL VDDHD VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] 
+ X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] 
+ XM[5] XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] 
+ YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I RTSEL[0]:I RTSEL[1]:I 
*.PININFO TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I 
*.PININFO X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I XM[0]:I XM[1]:I 
*.PININFO XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I Y[0]:I 
*.PININFO Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O 
*.PININFO BIST2IO:O BLEQ:O BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O 
*.PININFO DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O 
*.PININFO DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O 
*.PININFO DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O DEC_X2[5]:O 
*.PININFO DEC_X2[6]:O DEC_X2[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O 
*.PININFO DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O PD_BUF:O RE:O SAE:O 
*.PININFO VHI:O VLO:O WE:O YL[0]:O YL[1]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B
XCNT AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] 
+ DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] 
+ DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] 
+ DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] DEC_X2[5] 
+ DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] 
+ X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] 
+ XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3] 
+ S1AHSF400W40_CNT_CORE_884_BIST_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_884_BIST_M8M16_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_884_BIST_M8M16_SB AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB 
+ CEBM CKD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE 
+ TK TM TRKBL VDDHD VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] 
+ X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] 
+ XM[5] XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] 
+ YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I RTSEL[0]:I RTSEL[1]:I 
*.PININFO TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I 
*.PININFO X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I XM[0]:I XM[1]:I 
*.PININFO XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I Y[0]:I 
*.PININFO Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O 
*.PININFO BIST2IO:O BLEQ:O BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O 
*.PININFO DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O 
*.PININFO DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O 
*.PININFO DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O DEC_X2[5]:O 
*.PININFO DEC_X2[6]:O DEC_X2[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O 
*.PININFO DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O PD_BUF:O RE:O SAE:O 
*.PININFO VHI:O VLO:O WE:O YL[0]:O YL[1]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B
XCNT AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] 
+ DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] 
+ DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] 
+ DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] DEC_X2[5] 
+ DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] 
+ X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] 
+ XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3] 
+ S1AHSF400W40_CNT_CORE_884_BIST_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CDEC_M8_884_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CDEC_M8_884_SB BIST1B BIST2 BLEQ CEB CEBM CK1B CK2 CKD CKP CKPD CLK 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_Y[0] 
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN PD RE RSC 
+ VDDHD VDDI VSSI WE WEBXL WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] 
+ XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] Y[0] Y[1] Y[2] Y[3] YL[0] 
+ YL[1] YM[0] YM[1] YM[2] YM[3] AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7]
*.PININFO BIST1B:I BIST2:I CEB:I CEBM:I CKP:I CKPD:I CLK:I PD:I RSC:I WEBXL:I 
*.PININFO WEBXL1B:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I 
*.PININFO Y[0]:I Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I BLEQ:O 
*.PININFO CK1B:O CK2:O CKD:O DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O 
*.PININFO DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O DEC_X1[0]:O 
*.PININFO DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O DEC_X1[5]:O 
*.PININFO DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O DEC_X2[2]:O 
*.PININFO DEC_X2[3]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O 
*.PININFO DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O EN:O RE:O WE:O YL[0]:O YL[1]:O 
*.PININFO AX[0]:O AX[1]:O AX[2]:O AX[3]:O AX[4]:O AX[5]:O AX[6]:O AX[7]:O 
*.PININFO VDDHD:B VDDI:B VSSI:B
XIPDEC_X2<0> AXC[6] AXT[6] AXC[7] XC[0] XC[1] VDDHD VSSI S1AHSF400W40_DECB2_SB
XIPDEC_X2<1> AXC[6] AXT[6] AXT[7] XC[2] XC[3] VDDHD VSSI S1AHSF400W40_DECB2_SB
XIDEC_Y<0> NET0260 NET0260 DEC_Y[0] NET0260 NET0260 PD XY[0] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<1> NET0260 NET0260 DEC_Y[1] NET0260 NET0260 PD XY[1] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<2> NET0260 NET0260 DEC_Y[2] NET0260 NET0260 PD XY[2] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<3> NET0260 NET0260 DEC_Y[3] NET0260 NET0260 PD XY[3] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<4> NET0261 NET0261 DEC_Y[4] NET0261 NET0261 PD XY[4] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<5> NET0261 NET0261 DEC_Y[5] NET0261 NET0261 PD XY[5] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<6> NET0261 NET0261 DEC_Y[6] NET0261 NET0261 PD XY[6] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<7> NET0261 NET0261 DEC_Y[7] NET0261 NET0261 PD XY[7] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<0> NET0252 NET0252 DEC_X1[0] NET0252 NET0252 PD XB[0] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<1> NET0252 NET0252 DEC_X1[1] NET0252 NET0252 PD XB[1] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<2> NET0252 NET0252 DEC_X1[2] NET0252 NET0252 PD XB[2] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<3> NET0252 NET0252 DEC_X1[3] NET0252 NET0252 PD XB[3] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<4> NET0252 NET0252 DEC_X1[4] NET0252 NET0252 PD XB[4] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<5> NET0252 NET0252 DEC_X1[5] NET0252 NET0252 PD XB[5] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<6> NET0252 NET0252 DEC_X1[6] NET0252 NET0252 PD XB[6] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<7> NET0252 NET0252 DEC_X1[7] NET0252 NET0252 PD XB[7] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<0> NET0251 NET0251 DEC_X0[0] NET0251 NET0251 PD XA[0] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<1> NET0251 NET0251 DEC_X0[1] NET0251 NET0251 PD XA[1] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<2> NET0251 NET0251 DEC_X0[2] NET0251 NET0251 PD XA[2] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<3> NET0251 NET0251 DEC_X0[3] NET0251 NET0251 PD XA[3] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<4> NET0251 NET0251 DEC_X0[4] NET0251 NET0251 PD XA[4] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<5> NET0251 NET0251 DEC_X0[5] NET0251 NET0251 PD XA[5] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<6> NET0251 NET0251 DEC_X0[6] NET0251 NET0251 PD XA[6] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<7> NET0251 NET0251 DEC_X0[7] NET0251 NET0251 PD XA[7] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XDECB1_BLEQ BLEQ CKPD CLK_ENV ENC EN PD VDDHD VDDI VSSI S1AHSF400W40_DECB1_BLEQ_SB
XIPDEC_X0<0> AXC[0] AXT[0] AXC[1] AXT[1] AXC[2] XA[0] XA[1] XA[2] XA[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XIPDEC_X0<1> AXC[0] AXT[0] AXC[1] AXT[1] AXT[2] XA[4] XA[5] XA[6] XA[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XIPDEC_X1<0> AXC[3] AXT[3] AXC[4] AXT[4] AXC[5] XB[0] XB[1] XB[2] XB[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XIPDEC_X1<1> AXC[3] AXT[3] AXC[4] AXT[4] AXT[5] XB[4] XB[5] XB[6] XB[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XPREDEC_Y<0> AYC[0] AYT[0] AYC[1] AYT[1] AYC[2] XY[0] XY[1] XY[2] XY[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XPREDEC_Y<1> AYC[0] AYT[0] AYC[1] AYT[1] AYT[2] XY[4] XY[5] XY[6] XY[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XCKBUF CK1B CK2 CKPD CLK VDDHD VSSI S1AHSF400W40_CKBUF_SB
XABUF_Y<3> Y[3] YM[3] NET206 AYC[3] AYT[3] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<0> X[0] XM[0] AX[0] AXC[0] AXT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<1> X[1] XM[1] AX[1] AXC[1] AXT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<2> X[2] XM[2] AX[2] AXC[2] AXT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_Y<2> Y[2] YM[2] NET228 AYC[2] AYT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<6> X[6] XM[6] AX[6] AXC[6] AXT[6] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<7> X[7] XM[7] AX[7] AXC[7] AXT[7] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<3> X[3] XM[3] AX[3] AXC[3] AXT[3] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<4> X[4] XM[4] AX[4] AXC[4] AXT[4] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<5> X[5] XM[5] AX[5] AXC[5] AXT[5] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_Y<0> Y[0] YM[0] NET258[0] AYC[0] AYT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_Y<1> Y[1] YM[1] NET258[1] AYC[1] AYT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XCEBBUF BIST1B BIST2 CEB CEBM CK1B CK2 CKPD CLK CLK_ENV EN ENC RSC VDDHD VSSI 
+ S1AHSF400W40_ENBUFB_SB
XIDEC_REWE<0> CLK CLK_ENV RE EN ENC PD WEBXL VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_REWE<1> CLK CLK_ENV WE EN ENC PD WEBXL1B VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_CKD CLK CLK_ENV CKD EN ENC PD WEBXL1B VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_YL<0> CLK CLK_ENV YL[0] EN ENC PD AYC[3] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_YL<1> CLK CLK_ENV YL[1] EN ENC PD AYT[3] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<0> CLK CLK_ENV DEC_X2[0] EN ENC PD XC[0] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<1> CLK CLK_ENV DEC_X2[1] EN ENC PD XC[1] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<2> CLK CLK_ENV DEC_X2[2] EN ENC PD XC[2] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<3> CLK CLK_ENV DEC_X2[3] EN ENC PD XC[3] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    VHILO
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_VHILO VDDHD VHI VLO VSSI
*.PININFO VHI:O VLO:O VDDHD:B VSSI:B
MP0 Z2 Z2 VDDHD VDDHD PCH L=60N W=600N M=1
MP2 VHI Z1 VDDHD VDDHD PCH L=60N W=6U M=1
MP7 Z2 Z1 VDDHD VDDHD PCH L=60N W=600N M=1
MN1 VSSI Z2 VLO VSSI NCH L=60N W=6U M=2
MN0 VSSI Z1 Z1 VSSI NCH L=60N W=600N M=1
MN3 VSSI Z2 Z1 VSSI NCH L=60N W=600N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    COTH_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_COTH_SB AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKP 
+ CKPD CLK EN PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL VDDHD VDDI VHI 
+ VLO VSSI WEB WEBM WEBXL WEBXL1B WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] 
+ WTSEL[1] WTSEL[2]
*.PININFO AWT:I BIST:I CK1B:I CK2:I CLK:I EN:I PD:I PTSEL:I RTSEL[0]:I 
*.PININFO RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I AWT2:O 
*.PININFO BIST1B:O BIST2:O BIST2IO:O BLTRKWLDRV:O CKP:O CKPD:O PD_BUF:O RSC:O 
*.PININFO VHI:O VLO:O WEBXL:O WEBXL1B:O WLP_SAE:O WLP_SAEB:O TK:B TRKBL:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE_TK:B
MP1 VDDHD PD VDDI VDDI PCH L=60N W=3U M=9
MP0 VDDHD PD VDDI VDDI PCH L=60N W=3.8U M=16
XWEBBUF_SB BIST1B BIST2 CK1B CK2 VDDHD VSSI WEB WEBM WEBXL WEBXL1B S1AHSF400W40_WEBBUF_SB
XPDBUF_SB PD PD_BUF VDDI VSSI S1AHSF400W40_PDBUF_SB
XCKG CKP CLK EN RSC RSTCK TM VDDHD VSSI S1AHSF400W40_CKG_SB
XVHILO VDDHD VHI VLO VSSI S1AHSF400W40_VHILO
XRESETD BLTRKWLDRV CK2 CKP CKPD CKPDCLK WLP_SAEB RSTCK TK TRKBL VDDHD VSSI 
+ WEBXL WLP_SAE WLP_SAE_TK PTSEL RTSEL[0] RTSEL[1] WTSEL[0] WTSEL[1] WTSEL[2] 
+ S1AHSF400W40_RESETD_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_884_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_884_SB AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM CKD CLK 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] 
+ DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE TK TM 
+ TRKBL VDDHD VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] X[0] 
+ X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I RTSEL[0]:I RTSEL[1]:I 
*.PININFO TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I 
*.PININFO X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I XM[0]:I XM[1]:I 
*.PININFO XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I Y[0]:I 
*.PININFO Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O 
*.PININFO BIST2IO:O BLEQ:O BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O 
*.PININFO DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O 
*.PININFO DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O 
*.PININFO DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O DEC_X2[5]:O 
*.PININFO DEC_X2[6]:O DEC_X2[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O 
*.PININFO DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O PD_BUF:O RE:O SAE:O 
*.PININFO VHI:O VLO:O WE:O YL[0]:O YL[1]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B
XCDEC BIST1B BIST2 BLEQ CEB CEBM CK1B CK2 CKD CKP CKPD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN PD_BUF RE RSC VDDHD VDDI VSSI WE 
+ WEBXL WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] XM[0] XM[1] XM[2] 
+ XM[3] XM[4] XM[5] XM[6] XM[7] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] 
+ YM[2] YM[3] AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] S1AHSF400W40_CDEC_M8_884_SB
XCOTHERS AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKP CKPD CLK 
+ EN PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL VDDHD VDDI VHI VLO VSSI 
+ WEB WEBM WEBXL WEBXL1B SAE WLP_SAEB NET95 WTSEL[0] WTSEL[1] WTSEL[2] 
+ S1AHSF400W40_COTH_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_884_M4_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_884_M4_SB AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM CKD 
+ CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] 
+ DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE TK TM 
+ TRKBL VDDHD VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] X[0] 
+ X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I RTSEL[0]:I RTSEL[1]:I 
*.PININFO TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I 
*.PININFO X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I XM[0]:I XM[1]:I 
*.PININFO XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I Y[0]:I 
*.PININFO Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O 
*.PININFO BIST2IO:O BLEQ:O BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O 
*.PININFO DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O 
*.PININFO DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O 
*.PININFO DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O DEC_X2[5]:O 
*.PININFO DEC_X2[6]:O DEC_X2[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O 
*.PININFO DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O PD_BUF:O RE:O SAE:O 
*.PININFO VHI:O VLO:O WE:O YL[0]:O YL[1]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B
XCNT AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] 
+ DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] 
+ DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] 
+ DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] DEC_X2[5] 
+ DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] 
+ X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] 
+ XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3] 
+ S1AHSF400W40_CNT_CORE_884_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_884_M8M16_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_884_M8M16_SB AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM 
+ CKD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE 
+ TK TM TRKBL VDDHD VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] 
+ X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] 
+ XM[5] XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] 
+ YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I RTSEL[0]:I RTSEL[1]:I 
*.PININFO TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I 
*.PININFO X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I XM[0]:I XM[1]:I 
*.PININFO XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I Y[0]:I 
*.PININFO Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O 
*.PININFO BIST2IO:O BLEQ:O BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O 
*.PININFO DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O 
*.PININFO DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O 
*.PININFO DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O DEC_X2[5]:O 
*.PININFO DEC_X2[6]:O DEC_X2[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O 
*.PININFO DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O PD_BUF:O RE:O SAE:O 
*.PININFO VHI:O VLO:O WE:O YL[0]:O YL[1]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B
XCNT AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] 
+ DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] 
+ DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] 
+ DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] DEC_X2[5] 
+ DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] 
+ X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] 
+ XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3] 
+ S1AHSF400W40_CNT_CORE_884_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CDEC_M8_888_BIST_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CDEC_M8_888_BIST_SB BIST1B BIST2 BLEQ CEB CEBM CK1B CK2 CKD CKP CKPD 
+ CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] 
+ DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] EN PD RE RSC VDDHD VDDI VSSI WE WEBXL WEBXL1B 
+ X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] 
+ XM[5] XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] 
+ YM[3] AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8]
*.PININFO BIST1B:I BIST2:I CEB:I CEBM:I CKP:I CKPD:I CLK:I PD:I RSC:I WEBXL:I 
*.PININFO WEBXL1B:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I 
*.PININFO XM[7]:I XM[8]:I Y[0]:I Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I 
*.PININFO YM[3]:I BLEQ:O CK1B:O CK2:O CKD:O DEC_X0[0]:O DEC_X0[1]:O 
*.PININFO DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O 
*.PININFO DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O 
*.PININFO DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O DEC_X2[5]:O 
*.PININFO DEC_X2[6]:O DEC_X2[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O 
*.PININFO DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O EN:O RE:O WE:O YL[0]:O 
*.PININFO YL[1]:O AX[0]:O AX[1]:O AX[2]:O AX[3]:O AX[4]:O AX[5]:O AX[6]:O 
*.PININFO AX[7]:O AX[8]:O VDDHD:B VDDI:B VSSI:B
XCEBBUF BIST1B BIST2 CEB CEBM CK1B CK2 CKPD CLK CLK_ENV EN ENC RSC VDDHD VSSI 
+ S1AHSF400W40_ENBUFB_BIST_SB
XABUF_Y<3> Y[3] YM[3] NET161 AYC[3] AYT[3] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<6> X[6] XM[6] AX[6] AXC[6] AXT[6] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<7> X[7] XM[7] AX[7] AXC[7] AXT[7] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<8> X[8] XM[8] AX[8] AXC[8] AXT[8] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_Y<2> Y[2] YM[2] NET183 AYC[2] AYT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<3> X[3] XM[3] AX[3] AXC[3] AXT[3] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<4> X[4] XM[4] AX[4] AXC[4] AXT[4] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<5> X[5] XM[5] AX[5] AXC[5] AXT[5] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<0> X[0] XM[0] AX[0] AXC[0] AXT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<1> X[1] XM[1] AX[1] AXC[1] AXT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<2> X[2] XM[2] AX[2] AXC[2] AXT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_Y<0> Y[0] YM[0] NET213[0] AYC[0] AYT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_Y<1> Y[1] YM[1] NET213[1] AYC[1] AYT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XDECB1_BLEQ BLEQ CKPD CLK_ENV ENC EN PD VDDHD VDDI VSSI S1AHSF400W40_DECB1_BLEQ_SB
XIPDEC_X2<0> AXC[6] AXT[6] AXC[7] AXT[7] AXC[8] XC[0] XC[1] XC[2] XC[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XIPDEC_X2<1> AXC[6] AXT[6] AXC[7] AXT[7] AXT[8] XC[4] XC[5] XC[6] XC[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XIPDEC_X0<0> AXC[0] AXT[0] AXC[1] AXT[1] AXC[2] XA[0] XA[1] XA[2] XA[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XIPDEC_X0<1> AXC[0] AXT[0] AXC[1] AXT[1] AXT[2] XA[4] XA[5] XA[6] XA[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XPREDEC_Y<0> AYC[0] AYT[0] AYC[1] AYT[1] AYC[2] XY[0] XY[1] XY[2] XY[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XPREDEC_Y<1> AYC[0] AYT[0] AYC[1] AYT[1] AYT[2] XY[4] XY[5] XY[6] XY[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XIPDEC_X1<0> AXC[3] AXT[3] AXC[4] AXT[4] AXC[5] XB[0] XB[1] XB[2] XB[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XIPDEC_X1<1> AXC[3] AXT[3] AXC[4] AXT[4] AXT[5] XB[4] XB[5] XB[6] XB[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XCKBUF CK1B CK2 CKPD CLK VDDHD VSSI S1AHSF400W40_CKBUF_SB
XIDEC_Y<0> NET259 NET259 DEC_Y[0] NET259 NET259 PD XY[0] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<1> NET259 NET259 DEC_Y[1] NET259 NET259 PD XY[1] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<2> NET259 NET259 DEC_Y[2] NET259 NET259 PD XY[2] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<3> NET259 NET259 DEC_Y[3] NET259 NET259 PD XY[3] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<4> NET260 NET260 DEC_Y[4] NET260 NET260 PD XY[4] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<5> NET260 NET260 DEC_Y[5] NET260 NET260 PD XY[5] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<6> NET260 NET260 DEC_Y[6] NET260 NET260 PD XY[6] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<7> NET260 NET260 DEC_Y[7] NET260 NET260 PD XY[7] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<0> NET264 NET264 DEC_X1[0] NET264 NET264 PD XB[0] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<1> NET264 NET264 DEC_X1[1] NET264 NET264 PD XB[1] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<2> NET264 NET264 DEC_X1[2] NET264 NET264 PD XB[2] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<3> NET264 NET264 DEC_X1[3] NET264 NET264 PD XB[3] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<4> NET264 NET264 DEC_X1[4] NET264 NET264 PD XB[4] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<5> NET264 NET264 DEC_X1[5] NET264 NET264 PD XB[5] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<6> NET264 NET264 DEC_X1[6] NET264 NET264 PD XB[6] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<7> NET264 NET264 DEC_X1[7] NET264 NET264 PD XB[7] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<0> NET266 NET266 DEC_X0[0] NET266 NET266 PD XA[0] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<1> NET266 NET266 DEC_X0[1] NET266 NET266 PD XA[1] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<2> NET266 NET266 DEC_X0[2] NET266 NET266 PD XA[2] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<3> NET266 NET266 DEC_X0[3] NET266 NET266 PD XA[3] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<4> NET266 NET266 DEC_X0[4] NET266 NET266 PD XA[4] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<5> NET266 NET266 DEC_X0[5] NET266 NET266 PD XA[5] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<6> NET266 NET266 DEC_X0[6] NET266 NET266 PD XA[6] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<7> NET266 NET266 DEC_X0[7] NET266 NET266 PD XA[7] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_CKD CLK CLK_ENV CKD EN ENC PD WEBXL1B VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_REWE<0> CLK CLK_ENV RE EN ENC PD WEBXL VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_REWE<1> CLK CLK_ENV WE EN ENC PD WEBXL1B VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_YL<0> CLK CLK_ENV YL[0] EN ENC PD AYC[3] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_YL<1> CLK CLK_ENV YL[1] EN ENC PD AYT[3] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<0> CLK CLK_ENV DEC_X2[0] EN ENC PD XC[0] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<1> CLK CLK_ENV DEC_X2[1] EN ENC PD XC[1] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<2> CLK CLK_ENV DEC_X2[2] EN ENC PD XC[2] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<3> CLK CLK_ENV DEC_X2[3] EN ENC PD XC[3] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<4> CLK CLK_ENV DEC_X2[4] EN ENC PD XC[4] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<5> CLK CLK_ENV DEC_X2[5] EN ENC PD XC[5] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<6> CLK CLK_ENV DEC_X2[6] EN ENC PD XC[6] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<7> CLK CLK_ENV DEC_X2[7] EN ENC PD XC[7] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_888_BIST_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_888_BIST_SB AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM 
+ CKD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE 
+ TK TM TRKBL VDDHD VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] 
+ X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] 
+ XM[5] XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] 
+ YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I RTSEL[0]:I RTSEL[1]:I 
*.PININFO TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I 
*.PININFO X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I XM[0]:I XM[1]:I 
*.PININFO XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I Y[0]:I 
*.PININFO Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O 
*.PININFO BIST2IO:O BLEQ:O BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O 
*.PININFO DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O 
*.PININFO DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O 
*.PININFO DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O DEC_X2[5]:O 
*.PININFO DEC_X2[6]:O DEC_X2[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O 
*.PININFO DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O PD_BUF:O RE:O SAE:O 
*.PININFO VHI:O VLO:O WE:O YL[0]:O YL[1]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B
XCOTHERS AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKP CKPD CLK 
+ EN PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL VDDHD VDDI VHI VLO VSSI 
+ WEB WEBM WEBXL WEBXL1B SAE WLP_SAEB NET95 WTSEL[0] WTSEL[1] WTSEL[2] 
+ S1AHSF400W40_COTH_BIST_SB
XCDEC BIST1B BIST2 BLEQ CEB CEBM CK1B CK2 CKD CKP CKPD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] DEC_X2[5] DEC_X2[6] 
+ DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] 
+ DEC_Y[7] EN PD_BUF RE RSC VDDHD VDDI VSSI WE WEBXL WEBXL1B X[0] X[1] X[2] 
+ X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] 
+ XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3] AX[0] 
+ AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8] S1AHSF400W40_CDEC_M8_888_BIST_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_888_BIST_M4_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_888_BIST_M4_SB AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM 
+ CKD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE 
+ TK TM TRKBL VDDHD VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] 
+ X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] 
+ XM[5] XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] 
+ YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I RTSEL[0]:I RTSEL[1]:I 
*.PININFO TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I 
*.PININFO X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I XM[0]:I XM[1]:I 
*.PININFO XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I Y[0]:I 
*.PININFO Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O 
*.PININFO BIST2IO:O BLEQ:O BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O 
*.PININFO DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O 
*.PININFO DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O 
*.PININFO DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O DEC_X2[5]:O 
*.PININFO DEC_X2[6]:O DEC_X2[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O 
*.PININFO DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O PD_BUF:O RE:O SAE:O 
*.PININFO VHI:O VLO:O WE:O YL[0]:O YL[1]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B
XCNT AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] 
+ DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] 
+ DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] 
+ DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] DEC_X2[5] 
+ DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] 
+ X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] 
+ XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3] 
+ S1AHSF400W40_CNT_CORE_888_BIST_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_888_BIST_M8M16_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_888_BIST_M8M16_SB AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB 
+ CEBM CKD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE 
+ TK TM TRKBL VDDHD VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] 
+ X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] 
+ XM[5] XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] 
+ YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I RTSEL[0]:I RTSEL[1]:I 
*.PININFO TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I 
*.PININFO X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I XM[0]:I XM[1]:I 
*.PININFO XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I Y[0]:I 
*.PININFO Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O 
*.PININFO BIST2IO:O BLEQ:O BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O 
*.PININFO DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O 
*.PININFO DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O 
*.PININFO DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O DEC_X2[5]:O 
*.PININFO DEC_X2[6]:O DEC_X2[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O 
*.PININFO DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O PD_BUF:O RE:O SAE:O 
*.PININFO VHI:O VLO:O WE:O YL[0]:O YL[1]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B
XCNT AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] 
+ DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] 
+ DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] 
+ DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] DEC_X2[5] 
+ DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] 
+ X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] 
+ XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3] 
+ S1AHSF400W40_CNT_CORE_888_BIST_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CDEC_M8_888_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CDEC_M8_888_SB BIST1B BIST2 BLEQ CEB CEBM CK1B CK2 CKD CKP CKPD CLK 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] 
+ DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] EN PD RE RSC VDDHD VDDI VSSI WE WEBXL WEBXL1B 
+ X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] 
+ XM[5] XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] 
+ YM[3] AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8]
*.PININFO BIST1B:I BIST2:I CEB:I CEBM:I CKP:I CKPD:I CLK:I PD:I RSC:I WEBXL:I 
*.PININFO WEBXL1B:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I 
*.PININFO XM[7]:I XM[8]:I Y[0]:I Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I 
*.PININFO YM[3]:I BLEQ:O CK1B:O CK2:O CKD:O DEC_X0[0]:O DEC_X0[1]:O 
*.PININFO DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O 
*.PININFO DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O 
*.PININFO DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O DEC_X2[5]:O 
*.PININFO DEC_X2[6]:O DEC_X2[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O 
*.PININFO DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O EN:O RE:O WE:O YL[0]:O 
*.PININFO YL[1]:O AX[0]:O AX[1]:O AX[2]:O AX[3]:O AX[4]:O AX[5]:O AX[6]:O 
*.PININFO AX[7]:O AX[8]:O VDDHD:B VDDI:B VSSI:B
XDECB1_BLEQ BLEQ CKPD CLK_ENV ENC EN PD VDDHD VDDI VSSI S1AHSF400W40_DECB1_BLEQ_SB
XIPDEC_X2<0> AXC[6] AXT[6] AXC[7] AXT[7] AXC[8] XC[0] XC[1] XC[2] XC[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XIPDEC_X2<1> AXC[6] AXT[6] AXC[7] AXT[7] AXT[8] XC[4] XC[5] XC[6] XC[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XIPDEC_X0<0> AXC[0] AXT[0] AXC[1] AXT[1] AXC[2] XA[0] XA[1] XA[2] XA[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XIPDEC_X0<1> AXC[0] AXT[0] AXC[1] AXT[1] AXT[2] XA[4] XA[5] XA[6] XA[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XPREDEC_Y<0> AYC[0] AYT[0] AYC[1] AYT[1] AYC[2] XY[0] XY[1] XY[2] XY[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XPREDEC_Y<1> AYC[0] AYT[0] AYC[1] AYT[1] AYT[2] XY[4] XY[5] XY[6] XY[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XIPDEC_X1<0> AXC[3] AXT[3] AXC[4] AXT[4] AXC[5] XB[0] XB[1] XB[2] XB[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XIPDEC_X1<1> AXC[3] AXT[3] AXC[4] AXT[4] AXT[5] XB[4] XB[5] XB[6] XB[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4_SB
XCKBUF CK1B CK2 CKPD CLK VDDHD VSSI S1AHSF400W40_CKBUF_SB
XIDEC_Y<0> NET259 NET259 DEC_Y[0] NET259 NET259 PD XY[0] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<1> NET259 NET259 DEC_Y[1] NET259 NET259 PD XY[1] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<2> NET259 NET259 DEC_Y[2] NET259 NET259 PD XY[2] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<3> NET259 NET259 DEC_Y[3] NET259 NET259 PD XY[3] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<4> NET260 NET260 DEC_Y[4] NET260 NET260 PD XY[4] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<5> NET260 NET260 DEC_Y[5] NET260 NET260 PD XY[5] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<6> NET260 NET260 DEC_Y[6] NET260 NET260 PD XY[6] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_Y<7> NET260 NET260 DEC_Y[7] NET260 NET260 PD XY[7] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<0> NET264 NET264 DEC_X1[0] NET264 NET264 PD XB[0] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<1> NET264 NET264 DEC_X1[1] NET264 NET264 PD XB[1] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<2> NET264 NET264 DEC_X1[2] NET264 NET264 PD XB[2] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<3> NET264 NET264 DEC_X1[3] NET264 NET264 PD XB[3] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<4> NET264 NET264 DEC_X1[4] NET264 NET264 PD XB[4] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<5> NET264 NET264 DEC_X1[5] NET264 NET264 PD XB[5] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<6> NET264 NET264 DEC_X1[6] NET264 NET264 PD XB[6] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X1<7> NET264 NET264 DEC_X1[7] NET264 NET264 PD XB[7] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<0> NET266 NET266 DEC_X0[0] NET266 NET266 PD XA[0] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<1> NET266 NET266 DEC_X0[1] NET266 NET266 PD XA[1] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<2> NET266 NET266 DEC_X0[2] NET266 NET266 PD XA[2] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<3> NET266 NET266 DEC_X0[3] NET266 NET266 PD XA[3] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<4> NET266 NET266 DEC_X0[4] NET266 NET266 PD XA[4] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<5> NET266 NET266 DEC_X0[5] NET266 NET266 PD XA[5] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<6> NET266 NET266 DEC_X0[6] NET266 NET266 PD XA[6] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XIDEC_X0<7> NET266 NET266 DEC_X0[7] NET266 NET266 PD XA[7] VDDHD VSSI 
+ S1AHSF400W40_DECB1_X_SB
XABUF_Y<3> Y[3] YM[3] NET161 AYC[3] AYT[3] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<6> X[6] XM[6] AX[6] AXC[6] AXT[6] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<7> X[7] XM[7] AX[7] AXC[7] AXT[7] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<8> X[8] XM[8] AX[8] AXC[8] AXT[8] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_Y<2> Y[2] YM[2] NET183 AYC[2] AYT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<3> X[3] XM[3] AX[3] AXC[3] AXT[3] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<4> X[4] XM[4] AX[4] AXC[4] AXT[4] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<5> X[5] XM[5] AX[5] AXC[5] AXT[5] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<0> X[0] XM[0] AX[0] AXC[0] AXT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<1> X[1] XM[1] AX[1] AXC[1] AXT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<2> X[2] XM[2] AX[2] AXC[2] AXT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_Y<0> Y[0] YM[0] NET213[0] AYC[0] AYT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_Y<1> Y[1] YM[1] NET213[1] AYC[1] AYT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XCEBBUF BIST1B BIST2 CEB CEBM CK1B CK2 CKPD CLK CLK_ENV EN ENC RSC VDDHD VSSI 
+ S1AHSF400W40_ENBUFB_SB
XIDEC_CKD CLK CLK_ENV CKD EN ENC PD WEBXL1B VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_REWE<0> CLK CLK_ENV RE EN ENC PD WEBXL VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_REWE<1> CLK CLK_ENV WE EN ENC PD WEBXL1B VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_YL<0> CLK CLK_ENV YL[0] EN ENC PD AYC[3] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_YL<1> CLK CLK_ENV YL[1] EN ENC PD AYT[3] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<0> CLK CLK_ENV DEC_X2[0] EN ENC PD XC[0] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<1> CLK CLK_ENV DEC_X2[1] EN ENC PD XC[1] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<2> CLK CLK_ENV DEC_X2[2] EN ENC PD XC[2] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<3> CLK CLK_ENV DEC_X2[3] EN ENC PD XC[3] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<4> CLK CLK_ENV DEC_X2[4] EN ENC PD XC[4] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<5> CLK CLK_ENV DEC_X2[5] EN ENC PD XC[5] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<6> CLK CLK_ENV DEC_X2[6] EN ENC PD XC[6] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<7> CLK CLK_ENV DEC_X2[7] EN ENC PD XC[7] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_888_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_888_SB AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM CKD CLK 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] 
+ DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE TK TM 
+ TRKBL VDDHD VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] X[0] 
+ X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I RTSEL[0]:I RTSEL[1]:I 
*.PININFO TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I 
*.PININFO X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I XM[0]:I XM[1]:I 
*.PININFO XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I Y[0]:I 
*.PININFO Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O 
*.PININFO BIST2IO:O BLEQ:O BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O 
*.PININFO DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O 
*.PININFO DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O 
*.PININFO DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O DEC_X2[5]:O 
*.PININFO DEC_X2[6]:O DEC_X2[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O 
*.PININFO DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O PD_BUF:O RE:O SAE:O 
*.PININFO VHI:O VLO:O WE:O YL[0]:O YL[1]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B
XCDEC BIST1B BIST2 BLEQ CEB CEBM CK1B CK2 CKD CKP CKPD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] DEC_X2[5] DEC_X2[6] 
+ DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] 
+ DEC_Y[7] EN PD_BUF RE RSC VDDHD VDDI VSSI WE WEBXL WEBXL1B X[0] X[1] X[2] 
+ X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] 
+ XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3] AX[0] 
+ AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8] S1AHSF400W40_CDEC_M8_888_SB
XCOTHERS AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKP CKPD CLK 
+ EN PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL VDDHD VDDI VHI VLO VSSI 
+ WEB WEBM WEBXL WEBXL1B SAE WLP_SAEB NET95 WTSEL[0] WTSEL[1] WTSEL[2] 
+ S1AHSF400W40_COTH_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_888_M4_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_888_M4_SB AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM CKD 
+ CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] 
+ DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE TK TM 
+ TRKBL VDDHD VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] X[0] 
+ X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I RTSEL[0]:I RTSEL[1]:I 
*.PININFO TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I 
*.PININFO X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I XM[0]:I XM[1]:I 
*.PININFO XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I Y[0]:I 
*.PININFO Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O 
*.PININFO BIST2IO:O BLEQ:O BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O 
*.PININFO DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O 
*.PININFO DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O 
*.PININFO DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O DEC_X2[5]:O 
*.PININFO DEC_X2[6]:O DEC_X2[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O 
*.PININFO DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O PD_BUF:O RE:O SAE:O 
*.PININFO VHI:O VLO:O WE:O YL[0]:O YL[1]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B
XCNT AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] 
+ DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] 
+ DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] 
+ DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] DEC_X2[5] 
+ DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] 
+ X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] 
+ XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3] 
+ S1AHSF400W40_CNT_CORE_888_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_888_M8M16_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_888_M8M16_SB AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM 
+ CKD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE 
+ TK TM TRKBL VDDHD VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] 
+ X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] 
+ XM[5] XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] 
+ YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I RTSEL[0]:I RTSEL[1]:I 
*.PININFO TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I 
*.PININFO X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I XM[0]:I XM[1]:I 
*.PININFO XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I Y[0]:I 
*.PININFO Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O 
*.PININFO BIST2IO:O BLEQ:O BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O 
*.PININFO DEC_X0[2]:O DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O 
*.PININFO DEC_X0[7]:O DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O 
*.PININFO DEC_X1[4]:O DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O DEC_X2[5]:O 
*.PININFO DEC_X2[6]:O DEC_X2[7]:O DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O 
*.PININFO DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O DEC_Y[7]:O PD_BUF:O RE:O SAE:O 
*.PININFO VHI:O VLO:O WE:O YL[0]:O YL[1]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B
XCNT AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] 
+ DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] 
+ DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] 
+ DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] DEC_X2[5] 
+ DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] 
+ X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] 
+ XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3] 
+ S1AHSF400W40_CNT_CORE_888_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_CNT_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_CNT_SIM AWT AWT2 BIST BIST2IO BLEQ BLTRKWLDRV CEB CEBM CKD CLK 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] 
+ DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] PD PD_BUF PTSEL RE RTSEL[0] RTSEL[1] SAE TK TM 
+ TRKBL VDDHD VDDI VHI VLO VSSI WE WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] X[0] 
+ X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL[0] YL[1] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I RTSEL[0]:I RTSEL[1]:I 
*.PININFO TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I 
*.PININFO X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I XM[0]:I XM[1]:I 
*.PININFO XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I Y[0]:I 
*.PININFO Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:B 
*.PININFO BIST2IO:B BLEQ:B BLTRKWLDRV:B CKD:B DEC_X0[0]:B DEC_X0[1]:B 
*.PININFO DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B 
*.PININFO DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B 
*.PININFO DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B 
*.PININFO DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B DEC_X2[4]:B DEC_X2[5]:B 
*.PININFO DEC_X2[6]:B DEC_X2[7]:B DEC_Y[0]:B DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B 
*.PININFO DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B DEC_Y[7]:B PD_BUF:B RE:B SAE:B TK:B 
*.PININFO TRKBL:B VDDHD:B VDDI:B VHI:B VLO:B VSSI:B WE:B YL[0]:B YL[1]:B
XI311 NET51 NET60 NET50 NET56 NET53 NET59 NET49 NET48 NET58 NET47 NET42[0] 
+ NET42[1] NET42[2] NET42[3] NET42[4] NET42[5] NET42[6] NET42[7] NET62[0] 
+ NET62[1] NET62[2] NET62[3] NET62[4] NET62[5] NET62[6] NET62[7] NET72[0] 
+ NET72[1] NET72[2] NET72[3] NET72[4] NET72[5] NET72[6] NET72[7] NET71[0] 
+ NET71[1] NET71[2] NET71[3] NET71[4] NET71[5] NET71[6] NET71[7] NET46 NET41 
+ NET73 NET67 NET76[0] NET76[1] NET75 NET54 NET45 NET55 NET40 NET65 NET52 
+ NET57 NET64 NET69 NET44 NET43 NET74[0] NET74[1] NET74[2] NET63[0] NET63[1] 
+ NET63[2] NET63[3] NET63[4] NET63[5] NET63[6] NET63[7] NET63[8] NET61[0] 
+ NET61[1] NET61[2] NET61[3] NET61[4] NET61[5] NET61[6] NET61[7] NET61[8] 
+ NET70[0] NET70[1] NET70[2] NET70[3] NET66[0] NET66[1] NET68[0] NET68[1] 
+ NET68[2] NET68[3] S1AHSF400W40_CNT_CORE_882_BIST_M4_SB
XI312 NET88 NET97 NET87 NET93 NET90 NET96 NET86 NET85 NET95 NET84 NET79[0] 
+ NET79[1] NET79[2] NET79[3] NET79[4] NET79[5] NET79[6] NET79[7] NET99[0] 
+ NET99[1] NET99[2] NET99[3] NET99[4] NET99[5] NET99[6] NET99[7] NET109[0] 
+ NET109[1] NET109[2] NET109[3] NET109[4] NET109[5] NET109[6] NET109[7] 
+ NET108[0] NET108[1] NET108[2] NET108[3] NET108[4] NET108[5] NET108[6] 
+ NET108[7] NET83 NET78 NET110 NET104 NET113[0] NET113[1] NET112 NET91 NET82 
+ NET92 NET77 NET102 NET89 NET94 NET101 NET106 NET81 NET80 NET111[0] NET111[1] 
+ NET111[2] NET100[0] NET100[1] NET100[2] NET100[3] NET100[4] NET100[5] 
+ NET100[6] NET100[7] NET100[8] NET98[0] NET98[1] NET98[2] NET98[3] NET98[4] 
+ NET98[5] NET98[6] NET98[7] NET98[8] NET107[0] NET107[1] NET107[2] NET107[3] 
+ NET103[0] NET103[1] NET105[0] NET105[1] NET105[2] NET105[3] 
+ S1AHSF400W40_CNT_CORE_882_BIST_M8M16_SB
XI313 NET125 NET134 NET124 NET130 NET127 NET133 NET123 NET122 NET132 NET121 
+ NET116[0] NET116[1] NET116[2] NET116[3] NET116[4] NET116[5] NET116[6] 
+ NET116[7] NET136[0] NET136[1] NET136[2] NET136[3] NET136[4] NET136[5] 
+ NET136[6] NET136[7] NET146[0] NET146[1] NET146[2] NET146[3] NET146[4] 
+ NET146[5] NET146[6] NET146[7] NET145[0] NET145[1] NET145[2] NET145[3] 
+ NET145[4] NET145[5] NET145[6] NET145[7] NET120 NET115 NET147 NET141 
+ NET150[0] NET150[1] NET149 NET128 NET119 NET129 NET114 NET139 NET126 NET131 
+ NET138 NET143 NET118 NET117 NET148[0] NET148[1] NET148[2] NET137[0] 
+ NET137[1] NET137[2] NET137[3] NET137[4] NET137[5] NET137[6] NET137[7] 
+ NET137[8] NET135[0] NET135[1] NET135[2] NET135[3] NET135[4] NET135[5] 
+ NET135[6] NET135[7] NET135[8] NET144[0] NET144[1] NET144[2] NET144[3] 
+ NET140[0] NET140[1] NET142[0] NET142[1] NET142[2] NET142[3] 
+ S1AHSF400W40_CNT_CORE_882_M4_SB
XI314 NET162 NET171 NET161 NET167 NET164 NET170 NET160 NET159 NET169 NET158 
+ NET153[0] NET153[1] NET153[2] NET153[3] NET153[4] NET153[5] NET153[6] 
+ NET153[7] NET173[0] NET173[1] NET173[2] NET173[3] NET173[4] NET173[5] 
+ NET173[6] NET173[7] NET183[0] NET183[1] NET183[2] NET183[3] NET183[4] 
+ NET183[5] NET183[6] NET183[7] NET182[0] NET182[1] NET182[2] NET182[3] 
+ NET182[4] NET182[5] NET182[6] NET182[7] NET157 NET152 NET184 NET178 
+ NET187[0] NET187[1] NET186 NET165 NET156 NET166 NET151 NET176 NET163 NET168 
+ NET175 NET180 NET155 NET154 NET185[0] NET185[1] NET185[2] NET174[0] 
+ NET174[1] NET174[2] NET174[3] NET174[4] NET174[5] NET174[6] NET174[7] 
+ NET174[8] NET172[0] NET172[1] NET172[2] NET172[3] NET172[4] NET172[5] 
+ NET172[6] NET172[7] NET172[8] NET181[0] NET181[1] NET181[2] NET181[3] 
+ NET177[0] NET177[1] NET179[0] NET179[1] NET179[2] NET179[3] 
+ S1AHSF400W40_CNT_CORE_882_M8M16_SB
XI315 NET199 NET208 NET198 NET204 NET201 NET207 NET197 NET196 NET206 NET195 
+ NET190[0] NET190[1] NET190[2] NET190[3] NET190[4] NET190[5] NET190[6] 
+ NET190[7] NET210[0] NET210[1] NET210[2] NET210[3] NET210[4] NET210[5] 
+ NET210[6] NET210[7] NET220[0] NET220[1] NET220[2] NET220[3] NET220[4] 
+ NET220[5] NET220[6] NET220[7] NET219[0] NET219[1] NET219[2] NET219[3] 
+ NET219[4] NET219[5] NET219[6] NET219[7] NET194 NET189 NET221 NET215 
+ NET224[0] NET224[1] NET223 NET202 NET193 NET203 NET188 NET213 NET200 NET205 
+ NET212 NET217 NET192 NET191 NET222[0] NET222[1] NET222[2] NET211[0] 
+ NET211[1] NET211[2] NET211[3] NET211[4] NET211[5] NET211[6] NET211[7] 
+ NET211[8] NET209[0] NET209[1] NET209[2] NET209[3] NET209[4] NET209[5] 
+ NET209[6] NET209[7] NET209[8] NET218[0] NET218[1] NET218[2] NET218[3] 
+ NET214[0] NET214[1] NET216[0] NET216[1] NET216[2] NET216[3] 
+ S1AHSF400W40_CNT_CORE_884_BIST_M4_SB
XI316 NET236 NET245 NET235 NET241 NET238 NET244 NET234 NET233 NET243 NET232 
+ NET227[0] NET227[1] NET227[2] NET227[3] NET227[4] NET227[5] NET227[6] 
+ NET227[7] NET247[0] NET247[1] NET247[2] NET247[3] NET247[4] NET247[5] 
+ NET247[6] NET247[7] NET257[0] NET257[1] NET257[2] NET257[3] NET257[4] 
+ NET257[5] NET257[6] NET257[7] NET256[0] NET256[1] NET256[2] NET256[3] 
+ NET256[4] NET256[5] NET256[6] NET256[7] NET231 NET226 NET258 NET252 
+ NET261[0] NET261[1] NET260 NET239 NET230 NET240 NET225 NET250 NET237 NET242 
+ NET249 NET254 NET229 NET228 NET259[0] NET259[1] NET259[2] NET248[0] 
+ NET248[1] NET248[2] NET248[3] NET248[4] NET248[5] NET248[6] NET248[7] 
+ NET248[8] NET246[0] NET246[1] NET246[2] NET246[3] NET246[4] NET246[5] 
+ NET246[6] NET246[7] NET246[8] NET255[0] NET255[1] NET255[2] NET255[3] 
+ NET251[0] NET251[1] NET253[0] NET253[1] NET253[2] NET253[3] 
+ S1AHSF400W40_CNT_CORE_884_BIST_M8M16_SB
XI317 NET273 NET282 NET272 NET278 NET275 NET281 NET271 NET270 NET280 NET269 
+ NET264[0] NET264[1] NET264[2] NET264[3] NET264[4] NET264[5] NET264[6] 
+ NET264[7] NET284[0] NET284[1] NET284[2] NET284[3] NET284[4] NET284[5] 
+ NET284[6] NET284[7] NET294[0] NET294[1] NET294[2] NET294[3] NET294[4] 
+ NET294[5] NET294[6] NET294[7] NET293[0] NET293[1] NET293[2] NET293[3] 
+ NET293[4] NET293[5] NET293[6] NET293[7] NET268 NET263 NET295 NET289 
+ NET298[0] NET298[1] NET297 NET276 NET267 NET277 NET262 NET287 NET274 NET279 
+ NET286 NET291 NET266 NET265 NET296[0] NET296[1] NET296[2] NET285[0] 
+ NET285[1] NET285[2] NET285[3] NET285[4] NET285[5] NET285[6] NET285[7] 
+ NET285[8] NET283[0] NET283[1] NET283[2] NET283[3] NET283[4] NET283[5] 
+ NET283[6] NET283[7] NET283[8] NET292[0] NET292[1] NET292[2] NET292[3] 
+ NET288[0] NET288[1] NET290[0] NET290[1] NET290[2] NET290[3] 
+ S1AHSF400W40_CNT_CORE_884_M4_SB
XI318 NET310 NET319 NET309 NET315 NET312 NET318 NET308 NET307 NET317 NET306 
+ NET301[0] NET301[1] NET301[2] NET301[3] NET301[4] NET301[5] NET301[6] 
+ NET301[7] NET321[0] NET321[1] NET321[2] NET321[3] NET321[4] NET321[5] 
+ NET321[6] NET321[7] NET331[0] NET331[1] NET331[2] NET331[3] NET331[4] 
+ NET331[5] NET331[6] NET331[7] NET330[0] NET330[1] NET330[2] NET330[3] 
+ NET330[4] NET330[5] NET330[6] NET330[7] NET305 NET300 NET332 NET326 
+ NET335[0] NET335[1] NET334 NET313 NET304 NET314 NET299 NET324 NET311 NET316 
+ NET323 NET328 NET303 NET302 NET333[0] NET333[1] NET333[2] NET322[0] 
+ NET322[1] NET322[2] NET322[3] NET322[4] NET322[5] NET322[6] NET322[7] 
+ NET322[8] NET320[0] NET320[1] NET320[2] NET320[3] NET320[4] NET320[5] 
+ NET320[6] NET320[7] NET320[8] NET329[0] NET329[1] NET329[2] NET329[3] 
+ NET325[0] NET325[1] NET327[0] NET327[1] NET327[2] NET327[3] 
+ S1AHSF400W40_CNT_CORE_884_M8M16_SB
XI319 NET347 NET356 NET346 NET352 NET349 NET355 NET345 NET344 NET354 NET343 
+ NET338[0] NET338[1] NET338[2] NET338[3] NET338[4] NET338[5] NET338[6] 
+ NET338[7] NET358[0] NET358[1] NET358[2] NET358[3] NET358[4] NET358[5] 
+ NET358[6] NET358[7] NET368[0] NET368[1] NET368[2] NET368[3] NET368[4] 
+ NET368[5] NET368[6] NET368[7] NET367[0] NET367[1] NET367[2] NET367[3] 
+ NET367[4] NET367[5] NET367[6] NET367[7] NET342 NET337 NET369 NET363 
+ NET372[0] NET372[1] NET371 NET350 NET341 NET351 NET336 NET361 NET348 NET353 
+ NET360 NET365 NET340 NET339 NET370[0] NET370[1] NET370[2] NET359[0] 
+ NET359[1] NET359[2] NET359[3] NET359[4] NET359[5] NET359[6] NET359[7] 
+ NET359[8] NET357[0] NET357[1] NET357[2] NET357[3] NET357[4] NET357[5] 
+ NET357[6] NET357[7] NET357[8] NET366[0] NET366[1] NET366[2] NET366[3] 
+ NET362[0] NET362[1] NET364[0] NET364[1] NET364[2] NET364[3] 
+ S1AHSF400W40_CNT_CORE_888_BIST_M4_SB
XI320 NET384 NET393 NET383 NET389 NET386 NET392 NET382 NET381 NET391 NET380 
+ NET375[0] NET375[1] NET375[2] NET375[3] NET375[4] NET375[5] NET375[6] 
+ NET375[7] NET395[0] NET395[1] NET395[2] NET395[3] NET395[4] NET395[5] 
+ NET395[6] NET395[7] NET405[0] NET405[1] NET405[2] NET405[3] NET405[4] 
+ NET405[5] NET405[6] NET405[7] NET404[0] NET404[1] NET404[2] NET404[3] 
+ NET404[4] NET404[5] NET404[6] NET404[7] NET379 NET374 NET406 NET400 
+ NET409[0] NET409[1] NET408 NET387 NET378 NET388 NET373 NET398 NET385 NET390 
+ NET397 NET402 NET377 NET376 NET407[0] NET407[1] NET407[2] NET396[0] 
+ NET396[1] NET396[2] NET396[3] NET396[4] NET396[5] NET396[6] NET396[7] 
+ NET396[8] NET394[0] NET394[1] NET394[2] NET394[3] NET394[4] NET394[5] 
+ NET394[6] NET394[7] NET394[8] NET403[0] NET403[1] NET403[2] NET403[3] 
+ NET399[0] NET399[1] NET401[0] NET401[1] NET401[2] NET401[3] 
+ S1AHSF400W40_CNT_CORE_888_BIST_M8M16_SB
XI321 NET421 NET430 NET420 NET426 NET423 NET429 NET419 NET418 NET428 NET417 
+ NET412[0] NET412[1] NET412[2] NET412[3] NET412[4] NET412[5] NET412[6] 
+ NET412[7] NET432[0] NET432[1] NET432[2] NET432[3] NET432[4] NET432[5] 
+ NET432[6] NET432[7] NET442[0] NET442[1] NET442[2] NET442[3] NET442[4] 
+ NET442[5] NET442[6] NET442[7] NET441[0] NET441[1] NET441[2] NET441[3] 
+ NET441[4] NET441[5] NET441[6] NET441[7] NET416 NET411 NET443 NET437 
+ NET446[0] NET446[1] NET445 NET424 NET415 NET425 NET410 NET435 NET422 NET427 
+ NET434 NET439 NET414 NET413 NET444[0] NET444[1] NET444[2] NET433[0] 
+ NET433[1] NET433[2] NET433[3] NET433[4] NET433[5] NET433[6] NET433[7] 
+ NET433[8] NET431[0] NET431[1] NET431[2] NET431[3] NET431[4] NET431[5] 
+ NET431[6] NET431[7] NET431[8] NET440[0] NET440[1] NET440[2] NET440[3] 
+ NET436[0] NET436[1] NET438[0] NET438[1] NET438[2] NET438[3] 
+ S1AHSF400W40_CNT_CORE_888_M4_SB
XI322 NET458 NET467 NET457 NET463 NET460 NET466 NET456 NET455 NET465 NET454 
+ NET449[0] NET449[1] NET449[2] NET449[3] NET449[4] NET449[5] NET449[6] 
+ NET449[7] NET469[0] NET469[1] NET469[2] NET469[3] NET469[4] NET469[5] 
+ NET469[6] NET469[7] NET479[0] NET479[1] NET479[2] NET479[3] NET479[4] 
+ NET479[5] NET479[6] NET479[7] NET478[0] NET478[1] NET478[2] NET478[3] 
+ NET478[4] NET478[5] NET478[6] NET478[7] NET453 NET448 NET480 NET474 
+ NET483[0] NET483[1] NET482 NET461 NET452 NET462 NET447 NET472 NET459 NET464 
+ NET471 NET476 NET451 NET450 NET481[0] NET481[1] NET481[2] NET470[0] 
+ NET470[1] NET470[2] NET470[3] NET470[4] NET470[5] NET470[6] NET470[7] 
+ NET470[8] NET468[0] NET468[1] NET468[2] NET468[3] NET468[4] NET468[5] 
+ NET468[6] NET468[7] NET468[8] NET477[0] NET477[1] NET477[2] NET477[3] 
+ NET473[0] NET473[1] NET475[0] NET475[1] NET475[2] NET475[3] 
+ S1AHSF400W40_CNT_CORE_888_M8M16_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MCB_TKWL
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_TKWL BL BLB VDDI VSSI WL
*.PININFO BL:B BLB:B VDDI:B VSSI:B WL:B
MPCHPU1 FLOAT_MCB FLOAT_MC VDDI VDDI PCHPU_WISR L=0.065U W=0.080U M=1
MPCHPU0 VDDI FLOAT_MCB FLOAT_MC VDDI PCHPU_WISR L=0.065U W=0.080U M=1
MNCHPD1 BLB_IN FLOAT_MC VSSI VSSI NCHPD_WISR L=0.065U W=0.140U M=1
MNCHPD0 VSSI FLOAT_MCB BL_IN VSSI NCHPD_WISR L=0.065U W=0.140U M=1
MNCHPG1 BLB WL BLB_IN VSSI NCHPG_WISR L=0.075U W=0.090U M=1
MNCHPG0 BL_IN WL BL VSSI NCHPG_WISR L=0.075U W=0.090U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    TKWL_2X2
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TKWL_2X2 CVDDI VSSI WL_DUM WL_TK
*.PININFO CVDDI:B VSSI:B WL_DUM:B WL_TK:B
XTKWL_MCB_0 FLOAT_BL_L_T FLOAT_BLB_L CVDDI VSSI WL_TK S1AHSF400W40_MCB_TKWL
XTKDUM_MCB_1 FLOAT_BL_R_B FLOAT_BLB_R CVDDI VSSI WL_DUM S1AHSF400W40_MCB_TKWL
XTKWL_MCB_1 FLOAT_BL_R_T FLOAT_BLB_R CVDDI VSSI WL_TK S1AHSF400W40_MCB_TKWL
XTKDUM_MCB_0 FLOAT_BL_L_B FLOAT_BLB_L CVDDI VSSI WL_DUM S1AHSF400W40_MCB_TKWL
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    TKWL_LD_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TKWL_LD_SIM CVDDI TK_LT TK_RT VSSI WL_DUM_LT WL_DUM_RT WL_TK_LT 
+ WL_TK_RT
*.PININFO CVDDI:B TK_LT:B TK_RT:B VSSI:B WL_DUM_LT:B WL_DUM_RT:B WL_TK_LT:B 
*.PININFO WL_TK_RT:B
XI2 NET04 NET05 NET010 NET09 S1AHSF400W40_TKWL_2X2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    TKWL_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TKWL_SIM CVDDI TK_LT TK_RT VSSI WL_DUM_LT WL_DUM_RT WL_TK_LT WL_TK_RT
*.PININFO CVDDI:B TK_LT:B TK_RT:B VSSI:B WL_DUM_LT:B WL_DUM_RT:B WL_TK_LT:B 
*.PININFO WL_TK_RT:B
XTKWL_2X2 NET10 NET9 NET09 NET010 S1AHSF400W40_TKWL_2X2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SIM_SB1S
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SIM_SB1S AWT BIST BWEBM_LL BWEBM_LR BWEB_LL BWEB_LR CEB CEBM CLK DM_LL 
+ DM_LR D_LL D_LR PD PTSEL Q_LL Q_LR RTSEL[0] RTSEL[1] TM VDDI VSSI WEB WEBM 
+ WL_TK_ACT[0] WL_TK_ACT[1] WL_TK_ACT[2] WL_TK_ACT[3] WL_TK_ACT[4] 
+ WL_TK_ACT[5] WL_TK_ACT[6] WL_TK_ACT[7] WL_TK_ACT[8] WL_TK_ACT[9] 
+ WL_TK_ACT[10] WL_TK_ACT[11] WL_TK_ACT[12] WL_TK_ACT[13] WL_TK_ACT[14] 
+ WL_TK_ACT[15] WL_TK_ACT[16] WL_TK_ACT[17] WL_TK_ACT[18] WL_TK_ACT[19] 
+ WL_TK_ACT[20] WL_TK_ACT[21] WL_TK_ACT[22] WL_TK_ACT[23] WL_TK_ACT[24] 
+ WL_TK_ACT[25] WL_TK_ACT[26] WL_TK_ACT[27] WL_TK_ACT[28] WL_TK_ACT[29] 
+ WL_TK_ACT[30] WL_TK_ACT[31] WL_TK_ACT[32] WL_TK_ACT[33] WL_TK_ACT[34] 
+ WL_TK_ACT[35] WL_TK_ACT[36] WL_TK_ACT[37] WL_TK_ACT[38] WL_TK_ACT[39] 
+ WL_TK_ACT[40] WL_TK_ACT[41] WL_TK_ACT[42] WL_TK_ACT[43] WL_TK_ACT[44] 
+ WL_TK_ACT[45] WL_TK_ACT[46] WL_TK_ACT[47] WL_TK_ACT[48] WL_TK_ACT[49] 
+ WL_TK_ACT[50] WL_TK_ACT[51] WL_TK_ACT[52] WL_TK_ACT[53] WL_TK_ACT[54] 
+ WL_TK_ACT[55] WL_TK_ACT[56] WL_TK_ACT[57] WL_TK_ACT[58] WL_TK_ACT[59] 
+ WL_TK_ACT[60] WL_TK_ACT[61] WL_TK_ACT[62] WL_TK_ACT[63] WL_TK_ACT[64] 
+ WL_TK_ACT[65] WL_TK_ACT[66] WL_TK_ACT[67] WL_TK_ACT[68] WL_TK_ACT[69] 
+ WL_TK_ACT[70] WL_TK_ACT[71] WL_TK_ACT[72] WL_TK_ACT[73] WL_TK_ACT[74] 
+ WL_TK_ACT[75] WL_TK_ACT[76] WL_TK_ACT[77] WL_TK_ACT[78] WL_TK_ACT[79] 
+ WL_TK_ACT[80] WL_TK_ACT[81] WL_TK_ACT[82] WL_TK_ACT[83] WL_TK_ACT[84] 
+ WL_TK_ACT[85] WL_TK_ACT[86] WL_TK_ACT[87] WL_TK_ACT[88] WL_TK_ACT[89] 
+ WL_TK_ACT[90] WL_TK_ACT[91] WL_TK_ACT[92] WL_TK_ACT[93] WL_TK_ACT[94] 
+ WL_TK_ACT[95] WL_TK_ACT[96] WL_TK_ACT[97] WL_TK_ACT[98] WL_TK_ACT[99] 
+ WL_TK_ACT[100] WL_TK_ACT[101] WL_TK_ACT[102] WL_TK_ACT[103] WL_TK_ACT[104] 
+ WL_TK_ACT[105] WL_TK_ACT[106] WL_TK_ACT[107] WL_TK_ACT[108] WL_TK_ACT[109] 
+ WL_TK_ACT[110] WL_TK_ACT[111] WL_TK_ACT[112] WL_TK_ACT[113] WL_TK_ACT[114] 
+ WL_TK_ACT[115] WL_TK_ACT[116] WL_TK_ACT[117] WL_TK_ACT[118] WL_TK_ACT[119] 
+ WL_TK_ACT[120] WL_TK_ACT[121] WL_TK_ACT[122] WL_TK_ACT[123] WL_TK_ACT[124] 
+ WL_TK_ACT[125] WL_TK_ACT[126] WL_TK_ACT[127] WL_TK_ACT[128] WL_TK_ACT[129] 
+ WL_TK_ACT[130] WL_TK_ACT[131] WL_TK_ACT[132] WL_TK_ACT[133] WL_TK_ACT[134] 
+ WL_TK_ACT[135] WL_TK_ACT[136] WL_TK_ACT[137] WL_TK_ACT[138] WL_TK_ACT[139] 
+ WL_TK_ACT[140] WL_TK_ACT[141] WL_TK_ACT[142] WL_TK_ACT[143] WL_TK_ACT[144] 
+ WL_TK_ACT[145] WL_TK_ACT[146] WL_TK_ACT[147] WL_TK_ACT[148] WL_TK_ACT[149] 
+ WL_TK_ACT[150] WL_TK_ACT[151] WL_TK_ACT[152] WL_TK_ACT[153] WL_TK_ACT[154] 
+ WL_TK_ACT[155] WL_TK_ACT[156] WL_TK_ACT[157] WL_TK_ACT[158] WL_TK_ACT[159] 
+ WL_TK_ACT[160] WL_TK_ACT[161] WL_TK_ACT[162] WL_TK_ACT[163] WL_TK_ACT[164] 
+ WL_TK_ACT[165] WL_TK_ACT[166] WL_TK_ACT[167] WL_TK_ACT[168] WL_TK_ACT[169] 
+ WL_TK_ACT[170] WL_TK_ACT[171] WL_TK_ACT[172] WL_TK_ACT[173] WL_TK_ACT[174] 
+ WL_TK_ACT[175] WL_TK_ACT[176] WL_TK_ACT[177] WL_TK_ACT[178] WL_TK_ACT[179] 
+ WL_TK_ACT[180] WL_TK_ACT[181] WL_TK_ACT[182] WL_TK_ACT[183] WL_TK_ACT[184] 
+ WL_TK_ACT[185] WL_TK_ACT[186] WL_TK_ACT[187] WL_TK_ACT[188] WL_TK_ACT[189] 
+ WL_TK_ACT[190] WL_TK_ACT[191] WL_TK_ACT[192] WL_TK_ACT[193] WL_TK_ACT[194] 
+ WL_TK_ACT[195] WL_TK_ACT[196] WL_TK_ACT[197] WL_TK_ACT[198] WL_TK_ACT[199] 
+ WL_TK_ACT[200] WL_TK_ACT[201] WL_TK_ACT[202] WL_TK_ACT[203] WL_TK_ACT[204] 
+ WL_TK_ACT[205] WL_TK_ACT[206] WL_TK_ACT[207] WL_TK_ACT[208] WL_TK_ACT[209] 
+ WL_TK_ACT[210] WL_TK_ACT[211] WL_TK_ACT[212] WL_TK_ACT[213] WL_TK_ACT[214] 
+ WL_TK_ACT[215] WL_TK_ACT[216] WL_TK_ACT[217] WL_TK_ACT[218] WL_TK_ACT[219] 
+ WL_TK_ACT[220] WL_TK_ACT[221] WL_TK_ACT[222] WL_TK_ACT[223] WL_TK_ACT[224] 
+ WL_TK_ACT[225] WL_TK_ACT[226] WL_TK_ACT[227] WL_TK_ACT[228] WL_TK_ACT[229] 
+ WL_TK_ACT[230] WL_TK_ACT[231] WL_TK_ACT[232] WL_TK_ACT[233] WL_TK_ACT[234] 
+ WL_TK_ACT[235] WL_TK_ACT[236] WL_TK_ACT[237] WL_TK_ACT[238] WL_TK_ACT[239] 
+ WL_TK_ACT[240] WL_TK_ACT[241] WL_TK_ACT[242] WL_TK_ACT[243] WL_TK_ACT[244] 
+ WL_TK_ACT[245] WL_TK_ACT[246] WL_TK_ACT[247] WL_TK_ACT[248] WL_TK_ACT[249] 
+ WL_TK_ACT[250] WL_TK_ACT[251] WL_TK_ACT[252] WL_TK_ACT[253] WL_TK_ACT[254] 
+ WL_TK_ACT[255] WL_TK_ACT[256] WL_TK_ACT[257] WL_TK_ACT[258] WL_TK_ACT[259] 
+ WL_TK_ACT[260] WL_TK_ACT[261] WL_TK_ACT[262] WL_TK_ACT[263] WL_TK_ACT[264] 
+ WL_TK_ACT[265] WL_TK_ACT[266] WL_TK_ACT[267] WL_TK_ACT[268] WL_TK_ACT[269] 
+ WL_TK_ACT[270] WL_TK_ACT[271] WL_TK_ACT[272] WL_TK_ACT[273] WL_TK_ACT[274] 
+ WL_TK_ACT[275] WL_TK_ACT[276] WL_TK_ACT[277] WL_TK_ACT[278] WL_TK_ACT[279] 
+ WL_TK_ACT[280] WL_TK_ACT[281] WL_TK_ACT[282] WL_TK_ACT[283] WL_TK_ACT[284] 
+ WL_TK_ACT[285] WL_TK_ACT[286] WL_TK_ACT[287] WL_TK_ACT[288] WL_TK_ACT[289] 
+ WL_TK_ACT[290] WL_TK_ACT[291] WL_TK_ACT[292] WL_TK_ACT[293] WL_TK_ACT[294] 
+ WL_TK_ACT[295] WL_TK_ACT[296] WL_TK_ACT[297] WL_TK_ACT[298] WL_TK_ACT[299] 
+ WL_TK_ACT[300] WL_TK_ACT[301] WL_TK_ACT[302] WL_TK_ACT[303] WL_TK_ACT[304] 
+ WL_TK_ACT[305] WL_TK_ACT[306] WL_TK_ACT[307] WL_TK_ACT[308] WL_TK_ACT[309] 
+ WL_TK_ACT[310] WL_TK_ACT[311] WL_TK_ACT[312] WL_TK_ACT[313] WL_TK_ACT[314] 
+ WL_TK_ACT[315] WL_TK_ACT[316] WL_TK_ACT[317] WL_TK_ACT[318] WL_TK_ACT[319] 
+ WL_TK_ACT[320] WL_TK_ACT[321] WL_TK_ACT[322] WL_TK_ACT[323] WL_TK_ACT[324] 
+ WL_TK_ACT[325] WL_TK_ACT[326] WL_TK_ACT[327] WL_TK_ACT[328] WL_TK_ACT[329] 
+ WL_TK_ACT[330] WL_TK_ACT[331] WL_TK_ACT[332] WL_TK_ACT[333] WL_TK_ACT[334] 
+ WL_TK_ACT[335] WL_TK_ACT[336] WL_TK_ACT[337] WL_TK_ACT[338] WL_TK_ACT[339] 
+ WL_TK_ACT[340] WL_TK_ACT[341] WL_TK_ACT[342] WL_TK_ACT[343] WL_TK_ACT[344] 
+ WL_TK_ACT[345] WL_TK_ACT[346] WL_TK_ACT[347] WL_TK_ACT[348] WL_TK_ACT[349] 
+ WL_TK_ACT[350] WL_TK_ACT[351] WL_TK_ACT[352] WL_TK_ACT[353] WL_TK_ACT[354] 
+ WL_TK_ACT[355] WL_TK_ACT[356] WL_TK_ACT[357] WL_TK_ACT[358] WL_TK_ACT[359] 
+ WL_TK_ACT[360] WL_TK_ACT[361] WL_TK_ACT[362] WL_TK_ACT[363] WL_TK_ACT[364] 
+ WL_TK_ACT[365] WL_TK_ACT[366] WL_TK_ACT[367] WL_TK_ACT[368] WL_TK_ACT[369] 
+ WL_TK_ACT[370] WL_TK_ACT[371] WL_TK_ACT[372] WL_TK_ACT[373] WL_TK_ACT[374] 
+ WL_TK_ACT[375] WL_TK_ACT[376] WL_TK_ACT[377] WL_TK_ACT[378] WL_TK_ACT[379] 
+ WL_TK_ACT[380] WL_TK_ACT[381] WL_TK_ACT[382] WL_TK_ACT[383] WL_TK_ACT[384] 
+ WL_TK_ACT[385] WL_TK_ACT[386] WL_TK_ACT[387] WL_TK_ACT[388] WL_TK_ACT[389] 
+ WL_TK_ACT[390] WL_TK_ACT[391] WL_TK_ACT[392] WL_TK_ACT[393] WL_TK_ACT[394] 
+ WL_TK_ACT[395] WL_TK_ACT[396] WL_TK_ACT[397] WL_TK_ACT[398] WL_TK_ACT[399] 
+ WL_TK_ACT[400] WL_TK_ACT[401] WL_TK_ACT[402] WL_TK_ACT[403] WL_TK_ACT[404] 
+ WL_TK_ACT[405] WL_TK_ACT[406] WL_TK_ACT[407] WL_TK_ACT[408] WL_TK_ACT[409] 
+ WL_TK_ACT[410] WL_TK_ACT[411] WL_TK_ACT[412] WL_TK_ACT[413] WL_TK_ACT[414] 
+ WL_TK_ACT[415] WL_TK_ACT[416] WL_TK_ACT[417] WL_TK_ACT[418] WL_TK_ACT[419] 
+ WL_TK_ACT[420] WL_TK_ACT[421] WL_TK_ACT[422] WL_TK_ACT[423] WL_TK_ACT[424] 
+ WL_TK_ACT[425] WL_TK_ACT[426] WL_TK_ACT[427] WL_TK_ACT[428] WL_TK_ACT[429] 
+ WL_TK_ACT[430] WL_TK_ACT[431] WL_TK_ACT[432] WL_TK_ACT[433] WL_TK_ACT[434] 
+ WL_TK_ACT[435] WL_TK_ACT[436] WL_TK_ACT[437] WL_TK_ACT[438] WL_TK_ACT[439] 
+ WL_TK_ACT[440] WL_TK_ACT[441] WL_TK_ACT[442] WL_TK_ACT[443] WL_TK_ACT[444] 
+ WL_TK_ACT[445] WL_TK_ACT[446] WL_TK_ACT[447] WL_TK_ACT[448] WL_TK_ACT[449] 
+ WL_TK_ACT[450] WL_TK_ACT[451] WL_TK_ACT[452] WL_TK_ACT[453] WL_TK_ACT[454] 
+ WL_TK_ACT[455] WL_TK_ACT[456] WL_TK_ACT[457] WL_TK_ACT[458] WL_TK_ACT[459] 
+ WL_TK_ACT[460] WL_TK_ACT[461] WL_TK_ACT[462] WL_TK_ACT[463] WL_TK_ACT[464] 
+ WL_TK_ACT[465] WL_TK_ACT[466] WL_TK_ACT[467] WL_TK_ACT[468] WL_TK_ACT[469] 
+ WL_TK_ACT[470] WL_TK_ACT[471] WL_TK_ACT[472] WL_TK_ACT[473] WL_TK_ACT[474] 
+ WL_TK_ACT[475] WL_TK_ACT[476] WL_TK_ACT[477] WL_TK_ACT[478] WL_TK_ACT[479] 
+ WL_TK_ACT[480] WL_TK_ACT[481] WL_TK_ACT[482] WL_TK_ACT[483] WL_TK_ACT[484] 
+ WL_TK_ACT[485] WL_TK_ACT[486] WL_TK_ACT[487] WL_TK_ACT[488] WL_TK_ACT[489] 
+ WL_TK_ACT[490] WL_TK_ACT[491] WL_TK_ACT[492] WL_TK_ACT[493] WL_TK_ACT[494] 
+ WL_TK_ACT[495] WL_TK_ACT[496] WL_TK_ACT[497] WL_TK_ACT[498] WL_TK_ACT[499] 
+ WL_TK_ACT[500] WL_TK_ACT[501] WL_TK_ACT[502] WL_TK_ACT[503] WL_TK_ACT[504] 
+ WL_TK_ACT[505] WL_TK_ACT[506] WL_TK_ACT[507] WL_TK_ACT[508] WL_TK_ACT[509] 
+ WL_TK_ACT[510] WL_TK_ACT[511] WL_TK_LD WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] 
+ X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] 
+ XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I BWEBM_LL:I BWEBM_LR:I BWEB_LL:I BWEB_LR:I CEB:I CEBM:I 
*.PININFO CLK:I DM_LL:I DM_LR:I D_LL:I D_LR:I PD:I PTSEL:I RTSEL[0]:I 
*.PININFO RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I 
*.PININFO X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I XM[0]:I 
*.PININFO XM[1]:I XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I 
*.PININFO Y[0]:I Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I Q_LL:O 
*.PININFO Q_LR:O VDDI:B VSSI:B WL_TK_ACT[0]:B WL_TK_ACT[1]:B WL_TK_ACT[2]:B 
*.PININFO WL_TK_ACT[3]:B WL_TK_ACT[4]:B WL_TK_ACT[5]:B WL_TK_ACT[6]:B 
*.PININFO WL_TK_ACT[7]:B WL_TK_ACT[8]:B WL_TK_ACT[9]:B WL_TK_ACT[10]:B 
*.PININFO WL_TK_ACT[11]:B WL_TK_ACT[12]:B WL_TK_ACT[13]:B WL_TK_ACT[14]:B 
*.PININFO WL_TK_ACT[15]:B WL_TK_ACT[16]:B WL_TK_ACT[17]:B WL_TK_ACT[18]:B 
*.PININFO WL_TK_ACT[19]:B WL_TK_ACT[20]:B WL_TK_ACT[21]:B WL_TK_ACT[22]:B 
*.PININFO WL_TK_ACT[23]:B WL_TK_ACT[24]:B WL_TK_ACT[25]:B WL_TK_ACT[26]:B 
*.PININFO WL_TK_ACT[27]:B WL_TK_ACT[28]:B WL_TK_ACT[29]:B WL_TK_ACT[30]:B 
*.PININFO WL_TK_ACT[31]:B WL_TK_ACT[32]:B WL_TK_ACT[33]:B WL_TK_ACT[34]:B 
*.PININFO WL_TK_ACT[35]:B WL_TK_ACT[36]:B WL_TK_ACT[37]:B WL_TK_ACT[38]:B 
*.PININFO WL_TK_ACT[39]:B WL_TK_ACT[40]:B WL_TK_ACT[41]:B WL_TK_ACT[42]:B 
*.PININFO WL_TK_ACT[43]:B WL_TK_ACT[44]:B WL_TK_ACT[45]:B WL_TK_ACT[46]:B 
*.PININFO WL_TK_ACT[47]:B WL_TK_ACT[48]:B WL_TK_ACT[49]:B WL_TK_ACT[50]:B 
*.PININFO WL_TK_ACT[51]:B WL_TK_ACT[52]:B WL_TK_ACT[53]:B WL_TK_ACT[54]:B 
*.PININFO WL_TK_ACT[55]:B WL_TK_ACT[56]:B WL_TK_ACT[57]:B WL_TK_ACT[58]:B 
*.PININFO WL_TK_ACT[59]:B WL_TK_ACT[60]:B WL_TK_ACT[61]:B WL_TK_ACT[62]:B 
*.PININFO WL_TK_ACT[63]:B WL_TK_ACT[64]:B WL_TK_ACT[65]:B WL_TK_ACT[66]:B 
*.PININFO WL_TK_ACT[67]:B WL_TK_ACT[68]:B WL_TK_ACT[69]:B WL_TK_ACT[70]:B 
*.PININFO WL_TK_ACT[71]:B WL_TK_ACT[72]:B WL_TK_ACT[73]:B WL_TK_ACT[74]:B 
*.PININFO WL_TK_ACT[75]:B WL_TK_ACT[76]:B WL_TK_ACT[77]:B WL_TK_ACT[78]:B 
*.PININFO WL_TK_ACT[79]:B WL_TK_ACT[80]:B WL_TK_ACT[81]:B WL_TK_ACT[82]:B 
*.PININFO WL_TK_ACT[83]:B WL_TK_ACT[84]:B WL_TK_ACT[85]:B WL_TK_ACT[86]:B 
*.PININFO WL_TK_ACT[87]:B WL_TK_ACT[88]:B WL_TK_ACT[89]:B WL_TK_ACT[90]:B 
*.PININFO WL_TK_ACT[91]:B WL_TK_ACT[92]:B WL_TK_ACT[93]:B WL_TK_ACT[94]:B 
*.PININFO WL_TK_ACT[95]:B WL_TK_ACT[96]:B WL_TK_ACT[97]:B WL_TK_ACT[98]:B 
*.PININFO WL_TK_ACT[99]:B WL_TK_ACT[100]:B WL_TK_ACT[101]:B WL_TK_ACT[102]:B 
*.PININFO WL_TK_ACT[103]:B WL_TK_ACT[104]:B WL_TK_ACT[105]:B WL_TK_ACT[106]:B 
*.PININFO WL_TK_ACT[107]:B WL_TK_ACT[108]:B WL_TK_ACT[109]:B WL_TK_ACT[110]:B 
*.PININFO WL_TK_ACT[111]:B WL_TK_ACT[112]:B WL_TK_ACT[113]:B WL_TK_ACT[114]:B 
*.PININFO WL_TK_ACT[115]:B WL_TK_ACT[116]:B WL_TK_ACT[117]:B WL_TK_ACT[118]:B 
*.PININFO WL_TK_ACT[119]:B WL_TK_ACT[120]:B WL_TK_ACT[121]:B WL_TK_ACT[122]:B 
*.PININFO WL_TK_ACT[123]:B WL_TK_ACT[124]:B WL_TK_ACT[125]:B WL_TK_ACT[126]:B 
*.PININFO WL_TK_ACT[127]:B WL_TK_ACT[128]:B WL_TK_ACT[129]:B WL_TK_ACT[130]:B 
*.PININFO WL_TK_ACT[131]:B WL_TK_ACT[132]:B WL_TK_ACT[133]:B WL_TK_ACT[134]:B 
*.PININFO WL_TK_ACT[135]:B WL_TK_ACT[136]:B WL_TK_ACT[137]:B WL_TK_ACT[138]:B 
*.PININFO WL_TK_ACT[139]:B WL_TK_ACT[140]:B WL_TK_ACT[141]:B WL_TK_ACT[142]:B 
*.PININFO WL_TK_ACT[143]:B WL_TK_ACT[144]:B WL_TK_ACT[145]:B WL_TK_ACT[146]:B 
*.PININFO WL_TK_ACT[147]:B WL_TK_ACT[148]:B WL_TK_ACT[149]:B WL_TK_ACT[150]:B 
*.PININFO WL_TK_ACT[151]:B WL_TK_ACT[152]:B WL_TK_ACT[153]:B WL_TK_ACT[154]:B 
*.PININFO WL_TK_ACT[155]:B WL_TK_ACT[156]:B WL_TK_ACT[157]:B WL_TK_ACT[158]:B 
*.PININFO WL_TK_ACT[159]:B WL_TK_ACT[160]:B WL_TK_ACT[161]:B WL_TK_ACT[162]:B 
*.PININFO WL_TK_ACT[163]:B WL_TK_ACT[164]:B WL_TK_ACT[165]:B WL_TK_ACT[166]:B 
*.PININFO WL_TK_ACT[167]:B WL_TK_ACT[168]:B WL_TK_ACT[169]:B WL_TK_ACT[170]:B 
*.PININFO WL_TK_ACT[171]:B WL_TK_ACT[172]:B WL_TK_ACT[173]:B WL_TK_ACT[174]:B 
*.PININFO WL_TK_ACT[175]:B WL_TK_ACT[176]:B WL_TK_ACT[177]:B WL_TK_ACT[178]:B 
*.PININFO WL_TK_ACT[179]:B WL_TK_ACT[180]:B WL_TK_ACT[181]:B WL_TK_ACT[182]:B 
*.PININFO WL_TK_ACT[183]:B WL_TK_ACT[184]:B WL_TK_ACT[185]:B WL_TK_ACT[186]:B 
*.PININFO WL_TK_ACT[187]:B WL_TK_ACT[188]:B WL_TK_ACT[189]:B WL_TK_ACT[190]:B 
*.PININFO WL_TK_ACT[191]:B WL_TK_ACT[192]:B WL_TK_ACT[193]:B WL_TK_ACT[194]:B 
*.PININFO WL_TK_ACT[195]:B WL_TK_ACT[196]:B WL_TK_ACT[197]:B WL_TK_ACT[198]:B 
*.PININFO WL_TK_ACT[199]:B WL_TK_ACT[200]:B WL_TK_ACT[201]:B WL_TK_ACT[202]:B 
*.PININFO WL_TK_ACT[203]:B WL_TK_ACT[204]:B WL_TK_ACT[205]:B WL_TK_ACT[206]:B 
*.PININFO WL_TK_ACT[207]:B WL_TK_ACT[208]:B WL_TK_ACT[209]:B WL_TK_ACT[210]:B 
*.PININFO WL_TK_ACT[211]:B WL_TK_ACT[212]:B WL_TK_ACT[213]:B WL_TK_ACT[214]:B 
*.PININFO WL_TK_ACT[215]:B WL_TK_ACT[216]:B WL_TK_ACT[217]:B WL_TK_ACT[218]:B 
*.PININFO WL_TK_ACT[219]:B WL_TK_ACT[220]:B WL_TK_ACT[221]:B WL_TK_ACT[222]:B 
*.PININFO WL_TK_ACT[223]:B WL_TK_ACT[224]:B WL_TK_ACT[225]:B WL_TK_ACT[226]:B 
*.PININFO WL_TK_ACT[227]:B WL_TK_ACT[228]:B WL_TK_ACT[229]:B WL_TK_ACT[230]:B 
*.PININFO WL_TK_ACT[231]:B WL_TK_ACT[232]:B WL_TK_ACT[233]:B WL_TK_ACT[234]:B 
*.PININFO WL_TK_ACT[235]:B WL_TK_ACT[236]:B WL_TK_ACT[237]:B WL_TK_ACT[238]:B 
*.PININFO WL_TK_ACT[239]:B WL_TK_ACT[240]:B WL_TK_ACT[241]:B WL_TK_ACT[242]:B 
*.PININFO WL_TK_ACT[243]:B WL_TK_ACT[244]:B WL_TK_ACT[245]:B WL_TK_ACT[246]:B 
*.PININFO WL_TK_ACT[247]:B WL_TK_ACT[248]:B WL_TK_ACT[249]:B WL_TK_ACT[250]:B 
*.PININFO WL_TK_ACT[251]:B WL_TK_ACT[252]:B WL_TK_ACT[253]:B WL_TK_ACT[254]:B 
*.PININFO WL_TK_ACT[255]:B WL_TK_ACT[256]:B WL_TK_ACT[257]:B WL_TK_ACT[258]:B 
*.PININFO WL_TK_ACT[259]:B WL_TK_ACT[260]:B WL_TK_ACT[261]:B WL_TK_ACT[262]:B 
*.PININFO WL_TK_ACT[263]:B WL_TK_ACT[264]:B WL_TK_ACT[265]:B WL_TK_ACT[266]:B 
*.PININFO WL_TK_ACT[267]:B WL_TK_ACT[268]:B WL_TK_ACT[269]:B WL_TK_ACT[270]:B 
*.PININFO WL_TK_ACT[271]:B WL_TK_ACT[272]:B WL_TK_ACT[273]:B WL_TK_ACT[274]:B 
*.PININFO WL_TK_ACT[275]:B WL_TK_ACT[276]:B WL_TK_ACT[277]:B WL_TK_ACT[278]:B 
*.PININFO WL_TK_ACT[279]:B WL_TK_ACT[280]:B WL_TK_ACT[281]:B WL_TK_ACT[282]:B 
*.PININFO WL_TK_ACT[283]:B WL_TK_ACT[284]:B WL_TK_ACT[285]:B WL_TK_ACT[286]:B 
*.PININFO WL_TK_ACT[287]:B WL_TK_ACT[288]:B WL_TK_ACT[289]:B WL_TK_ACT[290]:B 
*.PININFO WL_TK_ACT[291]:B WL_TK_ACT[292]:B WL_TK_ACT[293]:B WL_TK_ACT[294]:B 
*.PININFO WL_TK_ACT[295]:B WL_TK_ACT[296]:B WL_TK_ACT[297]:B WL_TK_ACT[298]:B 
*.PININFO WL_TK_ACT[299]:B WL_TK_ACT[300]:B WL_TK_ACT[301]:B WL_TK_ACT[302]:B 
*.PININFO WL_TK_ACT[303]:B WL_TK_ACT[304]:B WL_TK_ACT[305]:B WL_TK_ACT[306]:B 
*.PININFO WL_TK_ACT[307]:B WL_TK_ACT[308]:B WL_TK_ACT[309]:B WL_TK_ACT[310]:B 
*.PININFO WL_TK_ACT[311]:B WL_TK_ACT[312]:B WL_TK_ACT[313]:B WL_TK_ACT[314]:B 
*.PININFO WL_TK_ACT[315]:B WL_TK_ACT[316]:B WL_TK_ACT[317]:B WL_TK_ACT[318]:B 
*.PININFO WL_TK_ACT[319]:B WL_TK_ACT[320]:B WL_TK_ACT[321]:B WL_TK_ACT[322]:B 
*.PININFO WL_TK_ACT[323]:B WL_TK_ACT[324]:B WL_TK_ACT[325]:B WL_TK_ACT[326]:B 
*.PININFO WL_TK_ACT[327]:B WL_TK_ACT[328]:B WL_TK_ACT[329]:B WL_TK_ACT[330]:B 
*.PININFO WL_TK_ACT[331]:B WL_TK_ACT[332]:B WL_TK_ACT[333]:B WL_TK_ACT[334]:B 
*.PININFO WL_TK_ACT[335]:B WL_TK_ACT[336]:B WL_TK_ACT[337]:B WL_TK_ACT[338]:B 
*.PININFO WL_TK_ACT[339]:B WL_TK_ACT[340]:B WL_TK_ACT[341]:B WL_TK_ACT[342]:B 
*.PININFO WL_TK_ACT[343]:B WL_TK_ACT[344]:B WL_TK_ACT[345]:B WL_TK_ACT[346]:B 
*.PININFO WL_TK_ACT[347]:B WL_TK_ACT[348]:B WL_TK_ACT[349]:B WL_TK_ACT[350]:B 
*.PININFO WL_TK_ACT[351]:B WL_TK_ACT[352]:B WL_TK_ACT[353]:B WL_TK_ACT[354]:B 
*.PININFO WL_TK_ACT[355]:B WL_TK_ACT[356]:B WL_TK_ACT[357]:B WL_TK_ACT[358]:B 
*.PININFO WL_TK_ACT[359]:B WL_TK_ACT[360]:B WL_TK_ACT[361]:B WL_TK_ACT[362]:B 
*.PININFO WL_TK_ACT[363]:B WL_TK_ACT[364]:B WL_TK_ACT[365]:B WL_TK_ACT[366]:B 
*.PININFO WL_TK_ACT[367]:B WL_TK_ACT[368]:B WL_TK_ACT[369]:B WL_TK_ACT[370]:B 
*.PININFO WL_TK_ACT[371]:B WL_TK_ACT[372]:B WL_TK_ACT[373]:B WL_TK_ACT[374]:B 
*.PININFO WL_TK_ACT[375]:B WL_TK_ACT[376]:B WL_TK_ACT[377]:B WL_TK_ACT[378]:B 
*.PININFO WL_TK_ACT[379]:B WL_TK_ACT[380]:B WL_TK_ACT[381]:B WL_TK_ACT[382]:B 
*.PININFO WL_TK_ACT[383]:B WL_TK_ACT[384]:B WL_TK_ACT[385]:B WL_TK_ACT[386]:B 
*.PININFO WL_TK_ACT[387]:B WL_TK_ACT[388]:B WL_TK_ACT[389]:B WL_TK_ACT[390]:B 
*.PININFO WL_TK_ACT[391]:B WL_TK_ACT[392]:B WL_TK_ACT[393]:B WL_TK_ACT[394]:B 
*.PININFO WL_TK_ACT[395]:B WL_TK_ACT[396]:B WL_TK_ACT[397]:B WL_TK_ACT[398]:B 
*.PININFO WL_TK_ACT[399]:B WL_TK_ACT[400]:B WL_TK_ACT[401]:B WL_TK_ACT[402]:B 
*.PININFO WL_TK_ACT[403]:B WL_TK_ACT[404]:B WL_TK_ACT[405]:B WL_TK_ACT[406]:B 
*.PININFO WL_TK_ACT[407]:B WL_TK_ACT[408]:B WL_TK_ACT[409]:B WL_TK_ACT[410]:B 
*.PININFO WL_TK_ACT[411]:B WL_TK_ACT[412]:B WL_TK_ACT[413]:B WL_TK_ACT[414]:B 
*.PININFO WL_TK_ACT[415]:B WL_TK_ACT[416]:B WL_TK_ACT[417]:B WL_TK_ACT[418]:B 
*.PININFO WL_TK_ACT[419]:B WL_TK_ACT[420]:B WL_TK_ACT[421]:B WL_TK_ACT[422]:B 
*.PININFO WL_TK_ACT[423]:B WL_TK_ACT[424]:B WL_TK_ACT[425]:B WL_TK_ACT[426]:B 
*.PININFO WL_TK_ACT[427]:B WL_TK_ACT[428]:B WL_TK_ACT[429]:B WL_TK_ACT[430]:B 
*.PININFO WL_TK_ACT[431]:B WL_TK_ACT[432]:B WL_TK_ACT[433]:B WL_TK_ACT[434]:B 
*.PININFO WL_TK_ACT[435]:B WL_TK_ACT[436]:B WL_TK_ACT[437]:B WL_TK_ACT[438]:B 
*.PININFO WL_TK_ACT[439]:B WL_TK_ACT[440]:B WL_TK_ACT[441]:B WL_TK_ACT[442]:B 
*.PININFO WL_TK_ACT[443]:B WL_TK_ACT[444]:B WL_TK_ACT[445]:B WL_TK_ACT[446]:B 
*.PININFO WL_TK_ACT[447]:B WL_TK_ACT[448]:B WL_TK_ACT[449]:B WL_TK_ACT[450]:B 
*.PININFO WL_TK_ACT[451]:B WL_TK_ACT[452]:B WL_TK_ACT[453]:B WL_TK_ACT[454]:B 
*.PININFO WL_TK_ACT[455]:B WL_TK_ACT[456]:B WL_TK_ACT[457]:B WL_TK_ACT[458]:B 
*.PININFO WL_TK_ACT[459]:B WL_TK_ACT[460]:B WL_TK_ACT[461]:B WL_TK_ACT[462]:B 
*.PININFO WL_TK_ACT[463]:B WL_TK_ACT[464]:B WL_TK_ACT[465]:B WL_TK_ACT[466]:B 
*.PININFO WL_TK_ACT[467]:B WL_TK_ACT[468]:B WL_TK_ACT[469]:B WL_TK_ACT[470]:B 
*.PININFO WL_TK_ACT[471]:B WL_TK_ACT[472]:B WL_TK_ACT[473]:B WL_TK_ACT[474]:B 
*.PININFO WL_TK_ACT[475]:B WL_TK_ACT[476]:B WL_TK_ACT[477]:B WL_TK_ACT[478]:B 
*.PININFO WL_TK_ACT[479]:B WL_TK_ACT[480]:B WL_TK_ACT[481]:B WL_TK_ACT[482]:B 
*.PININFO WL_TK_ACT[483]:B WL_TK_ACT[484]:B WL_TK_ACT[485]:B WL_TK_ACT[486]:B 
*.PININFO WL_TK_ACT[487]:B WL_TK_ACT[488]:B WL_TK_ACT[489]:B WL_TK_ACT[490]:B 
*.PININFO WL_TK_ACT[491]:B WL_TK_ACT[492]:B WL_TK_ACT[493]:B WL_TK_ACT[494]:B 
*.PININFO WL_TK_ACT[495]:B WL_TK_ACT[496]:B WL_TK_ACT[497]:B WL_TK_ACT[498]:B 
*.PININFO WL_TK_ACT[499]:B WL_TK_ACT[500]:B WL_TK_ACT[501]:B WL_TK_ACT[502]:B 
*.PININFO WL_TK_ACT[503]:B WL_TK_ACT[504]:B WL_TK_ACT[505]:B WL_TK_ACT[506]:B 
*.PININFO WL_TK_ACT[507]:B WL_TK_ACT[508]:B WL_TK_ACT[509]:B WL_TK_ACT[510]:B 
*.PININFO WL_TK_ACT[511]:B WL_TK_LD:B
XARR_WLLD_RD VDDI VDDHD VDDI VSSI WL_RD2[0] WL_RD2[1] WL_RD3[0] WL_RD3[1] 
+ S1AHSF400W40_SB_ARR_WLLD_SIM
XARR_WLLD_RU VDDI VDDHD VDDI VSSI WL_RU2[0] WL_RU2[1] WL_RU3[0] WL_RU3[1] 
+ S1AHSF400W40_SB_ARR_WLLD_SIM
XARR_WLLD_LD VDDI VDDHD VDDI VSSI WL_LD3[0] WL_LD3[1] WL_LD2[0] WL_LD2[1] 
+ S1AHSF400W40_SB_ARR_WLLD_SIM
XARR_WLLD_LU VDDI VDDHD VDDI VSSI WL_LU3[0] WL_LU3[1] WL_LU2[0] WL_LU2[1] 
+ S1AHSF400W40_SB_ARR_WLLD_SIM
XTKBL TRKBL BL_TK_TP VDDHD PD VDDHD VDDI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI WL_TK_ACT[0] 
+ WL_TK_ACT[1] WL_TK_ACT[2] WL_TK_ACT[3] WL_TK_ACT[4] WL_TK_ACT[5] 
+ WL_TK_ACT[6] WL_TK_ACT[7] WL_TK_ACT[8] WL_TK_ACT[9] WL_TK_ACT[10] 
+ WL_TK_ACT[11] WL_TK_ACT[12] WL_TK_ACT[13] WL_TK_ACT[14] WL_TK_ACT[15] 
+ WL_TK_ACT[16] WL_TK_ACT[17] WL_TK_ACT[18] WL_TK_ACT[19] WL_TK_ACT[20] 
+ WL_TK_ACT[21] WL_TK_ACT[22] WL_TK_ACT[23] WL_TK_ACT[24] WL_TK_ACT[25] 
+ WL_TK_ACT[26] WL_TK_ACT[27] WL_TK_ACT[28] WL_TK_ACT[29] WL_TK_ACT[30] 
+ WL_TK_ACT[31] WL_TK_ACT[32] WL_TK_ACT[33] WL_TK_ACT[34] WL_TK_ACT[35] 
+ WL_TK_ACT[36] WL_TK_ACT[37] WL_TK_ACT[38] WL_TK_ACT[39] WL_TK_ACT[40] 
+ WL_TK_ACT[41] WL_TK_ACT[42] WL_TK_ACT[43] WL_TK_ACT[44] WL_TK_ACT[45] 
+ WL_TK_ACT[46] WL_TK_ACT[47] WL_TK_ACT[48] WL_TK_ACT[49] WL_TK_ACT[50] 
+ WL_TK_ACT[51] WL_TK_ACT[52] WL_TK_ACT[53] WL_TK_ACT[54] WL_TK_ACT[55] 
+ WL_TK_ACT[56] WL_TK_ACT[57] WL_TK_ACT[58] WL_TK_ACT[59] WL_TK_ACT[60] 
+ WL_TK_ACT[61] WL_TK_ACT[62] WL_TK_ACT[63] WL_TK_ACT[64] WL_TK_ACT[65] 
+ WL_TK_ACT[66] WL_TK_ACT[67] WL_TK_ACT[68] WL_TK_ACT[69] WL_TK_ACT[70] 
+ WL_TK_ACT[71] WL_TK_ACT[72] WL_TK_ACT[73] WL_TK_ACT[74] WL_TK_ACT[75] 
+ WL_TK_ACT[76] WL_TK_ACT[77] WL_TK_ACT[78] WL_TK_ACT[79] WL_TK_ACT[80] 
+ WL_TK_ACT[81] WL_TK_ACT[82] WL_TK_ACT[83] WL_TK_ACT[84] WL_TK_ACT[85] 
+ WL_TK_ACT[86] WL_TK_ACT[87] WL_TK_ACT[88] WL_TK_ACT[89] WL_TK_ACT[90] 
+ WL_TK_ACT[91] WL_TK_ACT[92] WL_TK_ACT[93] WL_TK_ACT[94] WL_TK_ACT[95] 
+ WL_TK_ACT[96] WL_TK_ACT[97] WL_TK_ACT[98] WL_TK_ACT[99] WL_TK_ACT[100] 
+ WL_TK_ACT[101] WL_TK_ACT[102] WL_TK_ACT[103] WL_TK_ACT[104] WL_TK_ACT[105] 
+ WL_TK_ACT[106] WL_TK_ACT[107] WL_TK_ACT[108] WL_TK_ACT[109] WL_TK_ACT[110] 
+ WL_TK_ACT[111] WL_TK_ACT[112] WL_TK_ACT[113] WL_TK_ACT[114] WL_TK_ACT[115] 
+ WL_TK_ACT[116] WL_TK_ACT[117] WL_TK_ACT[118] WL_TK_ACT[119] WL_TK_ACT[120] 
+ WL_TK_ACT[121] WL_TK_ACT[122] WL_TK_ACT[123] WL_TK_ACT[124] WL_TK_ACT[125] 
+ WL_TK_ACT[126] WL_TK_ACT[127] WL_TK_ACT[128] WL_TK_ACT[129] WL_TK_ACT[130] 
+ WL_TK_ACT[131] WL_TK_ACT[132] WL_TK_ACT[133] WL_TK_ACT[134] WL_TK_ACT[135] 
+ WL_TK_ACT[136] WL_TK_ACT[137] WL_TK_ACT[138] WL_TK_ACT[139] WL_TK_ACT[140] 
+ WL_TK_ACT[141] WL_TK_ACT[142] WL_TK_ACT[143] WL_TK_ACT[144] WL_TK_ACT[145] 
+ WL_TK_ACT[146] WL_TK_ACT[147] WL_TK_ACT[148] WL_TK_ACT[149] WL_TK_ACT[150] 
+ WL_TK_ACT[151] WL_TK_ACT[152] WL_TK_ACT[153] WL_TK_ACT[154] WL_TK_ACT[155] 
+ WL_TK_ACT[156] WL_TK_ACT[157] WL_TK_ACT[158] WL_TK_ACT[159] WL_TK_ACT[160] 
+ WL_TK_ACT[161] WL_TK_ACT[162] WL_TK_ACT[163] WL_TK_ACT[164] WL_TK_ACT[165] 
+ WL_TK_ACT[166] WL_TK_ACT[167] WL_TK_ACT[168] WL_TK_ACT[169] WL_TK_ACT[170] 
+ WL_TK_ACT[171] WL_TK_ACT[172] WL_TK_ACT[173] WL_TK_ACT[174] WL_TK_ACT[175] 
+ WL_TK_ACT[176] WL_TK_ACT[177] WL_TK_ACT[178] WL_TK_ACT[179] WL_TK_ACT[180] 
+ WL_TK_ACT[181] WL_TK_ACT[182] WL_TK_ACT[183] WL_TK_ACT[184] WL_TK_ACT[185] 
+ WL_TK_ACT[186] WL_TK_ACT[187] WL_TK_ACT[188] WL_TK_ACT[189] WL_TK_ACT[190] 
+ WL_TK_ACT[191] WL_TK_ACT[192] WL_TK_ACT[193] WL_TK_ACT[194] WL_TK_ACT[195] 
+ WL_TK_ACT[196] WL_TK_ACT[197] WL_TK_ACT[198] WL_TK_ACT[199] WL_TK_ACT[200] 
+ WL_TK_ACT[201] WL_TK_ACT[202] WL_TK_ACT[203] WL_TK_ACT[204] WL_TK_ACT[205] 
+ WL_TK_ACT[206] WL_TK_ACT[207] WL_TK_ACT[208] WL_TK_ACT[209] WL_TK_ACT[210] 
+ WL_TK_ACT[211] WL_TK_ACT[212] WL_TK_ACT[213] WL_TK_ACT[214] WL_TK_ACT[215] 
+ WL_TK_ACT[216] WL_TK_ACT[217] WL_TK_ACT[218] WL_TK_ACT[219] WL_TK_ACT[220] 
+ WL_TK_ACT[221] WL_TK_ACT[222] WL_TK_ACT[223] WL_TK_ACT[224] WL_TK_ACT[225] 
+ WL_TK_ACT[226] WL_TK_ACT[227] WL_TK_ACT[228] WL_TK_ACT[229] WL_TK_ACT[230] 
+ WL_TK_ACT[231] WL_TK_ACT[232] WL_TK_ACT[233] WL_TK_ACT[234] WL_TK_ACT[235] 
+ WL_TK_ACT[236] WL_TK_ACT[237] WL_TK_ACT[238] WL_TK_ACT[239] WL_TK_ACT[240] 
+ WL_TK_ACT[241] WL_TK_ACT[242] WL_TK_ACT[243] WL_TK_ACT[244] WL_TK_ACT[245] 
+ WL_TK_ACT[246] WL_TK_ACT[247] WL_TK_ACT[248] WL_TK_ACT[249] WL_TK_ACT[250] 
+ WL_TK_ACT[251] WL_TK_ACT[252] WL_TK_ACT[253] WL_TK_ACT[254] WL_TK_ACT[255] 
+ WL_TK_ACT[256] WL_TK_ACT[257] WL_TK_ACT[258] WL_TK_ACT[259] WL_TK_ACT[260] 
+ WL_TK_ACT[261] WL_TK_ACT[262] WL_TK_ACT[263] WL_TK_ACT[264] WL_TK_ACT[265] 
+ WL_TK_ACT[266] WL_TK_ACT[267] WL_TK_ACT[268] WL_TK_ACT[269] WL_TK_ACT[270] 
+ WL_TK_ACT[271] WL_TK_ACT[272] WL_TK_ACT[273] WL_TK_ACT[274] WL_TK_ACT[275] 
+ WL_TK_ACT[276] WL_TK_ACT[277] WL_TK_ACT[278] WL_TK_ACT[279] WL_TK_ACT[280] 
+ WL_TK_ACT[281] WL_TK_ACT[282] WL_TK_ACT[283] WL_TK_ACT[284] WL_TK_ACT[285] 
+ WL_TK_ACT[286] WL_TK_ACT[287] WL_TK_ACT[288] WL_TK_ACT[289] WL_TK_ACT[290] 
+ WL_TK_ACT[291] WL_TK_ACT[292] WL_TK_ACT[293] WL_TK_ACT[294] WL_TK_ACT[295] 
+ WL_TK_ACT[296] WL_TK_ACT[297] WL_TK_ACT[298] WL_TK_ACT[299] WL_TK_ACT[300] 
+ WL_TK_ACT[301] WL_TK_ACT[302] WL_TK_ACT[303] WL_TK_ACT[304] WL_TK_ACT[305] 
+ WL_TK_ACT[306] WL_TK_ACT[307] WL_TK_ACT[308] WL_TK_ACT[309] WL_TK_ACT[310] 
+ WL_TK_ACT[311] WL_TK_ACT[312] WL_TK_ACT[313] WL_TK_ACT[314] WL_TK_ACT[315] 
+ WL_TK_ACT[316] WL_TK_ACT[317] WL_TK_ACT[318] WL_TK_ACT[319] WL_TK_ACT[320] 
+ WL_TK_ACT[321] WL_TK_ACT[322] WL_TK_ACT[323] WL_TK_ACT[324] WL_TK_ACT[325] 
+ WL_TK_ACT[326] WL_TK_ACT[327] WL_TK_ACT[328] WL_TK_ACT[329] WL_TK_ACT[330] 
+ WL_TK_ACT[331] WL_TK_ACT[332] WL_TK_ACT[333] WL_TK_ACT[334] WL_TK_ACT[335] 
+ WL_TK_ACT[336] WL_TK_ACT[337] WL_TK_ACT[338] WL_TK_ACT[339] WL_TK_ACT[340] 
+ WL_TK_ACT[341] WL_TK_ACT[342] WL_TK_ACT[343] WL_TK_ACT[344] WL_TK_ACT[345] 
+ WL_TK_ACT[346] WL_TK_ACT[347] WL_TK_ACT[348] WL_TK_ACT[349] WL_TK_ACT[350] 
+ WL_TK_ACT[351] WL_TK_ACT[352] WL_TK_ACT[353] WL_TK_ACT[354] WL_TK_ACT[355] 
+ WL_TK_ACT[356] WL_TK_ACT[357] WL_TK_ACT[358] WL_TK_ACT[359] WL_TK_ACT[360] 
+ WL_TK_ACT[361] WL_TK_ACT[362] WL_TK_ACT[363] WL_TK_ACT[364] WL_TK_ACT[365] 
+ WL_TK_ACT[366] WL_TK_ACT[367] WL_TK_ACT[368] WL_TK_ACT[369] WL_TK_ACT[370] 
+ WL_TK_ACT[371] WL_TK_ACT[372] WL_TK_ACT[373] WL_TK_ACT[374] WL_TK_ACT[375] 
+ WL_TK_ACT[376] WL_TK_ACT[377] WL_TK_ACT[378] WL_TK_ACT[379] WL_TK_ACT[380] 
+ WL_TK_ACT[381] WL_TK_ACT[382] WL_TK_ACT[383] WL_TK_ACT[384] WL_TK_ACT[385] 
+ WL_TK_ACT[386] WL_TK_ACT[387] WL_TK_ACT[388] WL_TK_ACT[389] WL_TK_ACT[390] 
+ WL_TK_ACT[391] WL_TK_ACT[392] WL_TK_ACT[393] WL_TK_ACT[394] WL_TK_ACT[395] 
+ WL_TK_ACT[396] WL_TK_ACT[397] WL_TK_ACT[398] WL_TK_ACT[399] WL_TK_ACT[400] 
+ WL_TK_ACT[401] WL_TK_ACT[402] WL_TK_ACT[403] WL_TK_ACT[404] WL_TK_ACT[405] 
+ WL_TK_ACT[406] WL_TK_ACT[407] WL_TK_ACT[408] WL_TK_ACT[409] WL_TK_ACT[410] 
+ WL_TK_ACT[411] WL_TK_ACT[412] WL_TK_ACT[413] WL_TK_ACT[414] WL_TK_ACT[415] 
+ WL_TK_ACT[416] WL_TK_ACT[417] WL_TK_ACT[418] WL_TK_ACT[419] WL_TK_ACT[420] 
+ WL_TK_ACT[421] WL_TK_ACT[422] WL_TK_ACT[423] WL_TK_ACT[424] WL_TK_ACT[425] 
+ WL_TK_ACT[426] WL_TK_ACT[427] WL_TK_ACT[428] WL_TK_ACT[429] WL_TK_ACT[430] 
+ WL_TK_ACT[431] WL_TK_ACT[432] WL_TK_ACT[433] WL_TK_ACT[434] WL_TK_ACT[435] 
+ WL_TK_ACT[436] WL_TK_ACT[437] WL_TK_ACT[438] WL_TK_ACT[439] WL_TK_ACT[440] 
+ WL_TK_ACT[441] WL_TK_ACT[442] WL_TK_ACT[443] WL_TK_ACT[444] WL_TK_ACT[445] 
+ WL_TK_ACT[446] WL_TK_ACT[447] WL_TK_ACT[448] WL_TK_ACT[449] WL_TK_ACT[450] 
+ WL_TK_ACT[451] WL_TK_ACT[452] WL_TK_ACT[453] WL_TK_ACT[454] WL_TK_ACT[455] 
+ WL_TK_ACT[456] WL_TK_ACT[457] WL_TK_ACT[458] WL_TK_ACT[459] WL_TK_ACT[460] 
+ WL_TK_ACT[461] WL_TK_ACT[462] WL_TK_ACT[463] WL_TK_ACT[464] WL_TK_ACT[465] 
+ WL_TK_ACT[466] WL_TK_ACT[467] WL_TK_ACT[468] WL_TK_ACT[469] WL_TK_ACT[470] 
+ WL_TK_ACT[471] WL_TK_ACT[472] WL_TK_ACT[473] WL_TK_ACT[474] WL_TK_ACT[475] 
+ WL_TK_ACT[476] WL_TK_ACT[477] WL_TK_ACT[478] WL_TK_ACT[479] WL_TK_ACT[480] 
+ WL_TK_ACT[481] WL_TK_ACT[482] WL_TK_ACT[483] WL_TK_ACT[484] WL_TK_ACT[485] 
+ WL_TK_ACT[486] WL_TK_ACT[487] WL_TK_ACT[488] WL_TK_ACT[489] WL_TK_ACT[490] 
+ WL_TK_ACT[491] WL_TK_ACT[492] WL_TK_ACT[493] WL_TK_ACT[494] WL_TK_ACT[495] 
+ WL_TK_ACT[496] WL_TK_ACT[497] WL_TK_ACT[498] WL_TK_ACT[499] WL_TK_ACT[500] 
+ WL_TK_ACT[501] WL_TK_ACT[502] WL_TK_ACT[503] WL_TK_ACT[504] WL_TK_ACT[505] 
+ WL_TK_ACT[506] WL_TK_ACT[507] WL_TK_ACT[508] WL_TK_ACT[509] WL_TK_ACT[510] 
+ WL_TK_ACT[511] TIEH_BT TIEL S1AHSF400W40_TKBL_SIM
XTRKPRE PD TRKBL WL_TK VDDHD VDDI VSSI TIEH_BT TIEL S1AHSF400W40_TRKPRE_SIM
XBK_WLDV_D DEC_X0_1[0] DEC_X0_1[1] DEC_X0_1[2] DEC_X0_1[3] DEC_X0_1[4] 
+ DEC_X0_1[5] DEC_X0_1[6] DEC_X0_1[7] DEC_X0_2[0] DEC_X0_2[1] DEC_X0_2[2] 
+ DEC_X0_2[3] DEC_X0_2[4] DEC_X0_2[5] DEC_X0_2[6] DEC_X0_2[7] DEC_X1_1[0] 
+ DEC_X1_1[1] DEC_X1_1[2] DEC_X1_1[3] DEC_X1_1[4] DEC_X1_1[5] DEC_X1_1[6] 
+ DEC_X1_1[7] DEC_X1_2[0] DEC_X1_2[1] DEC_X1_2[2] DEC_X1_2[3] DEC_X1_2[4] 
+ DEC_X1_2[5] DEC_X1_2[6] DEC_X1_2[7] DEC_X2_1[0] DEC_X2_1[1] DEC_X2_1[2] 
+ DEC_X2_1[3] DEC_X2_1[4] DEC_X2_1[5] DEC_X2_1[6] DEC_X2_1[7] DEC_X2_SHARE_2 
+ DEC_X2_2[0] DEC_X2_2[1] DEC_X2_2[2] DEC_X2_2[3] DEC_X2_2[4] DEC_X2_2[5] 
+ DEC_X2_2[6] DEC_X2_2[7] PD_BUF_L1 PD_BUF_2 VDDHD VDDI VSSI WL_LD1[0] 
+ WL_LD1[1] WL_RD1[0] WL_RD1[1] S1AHSF400W40_SB_WLDV_D_SIM
XBK_WLDV_U DEC_X0_3[0] DEC_X0_3[1] DEC_X0_3[2] DEC_X0_3[3] DEC_X0_3[4] 
+ DEC_X0_3[5] DEC_X0_3[6] DEC_X0_3[7] NET0132[0] NET0132[1] NET0132[2] 
+ NET0132[3] NET0132[4] NET0132[5] NET0132[6] NET0132[7] DEC_X1_3[0] 
+ DEC_X1_3[1] DEC_X1_3[2] DEC_X1_3[3] DEC_X1_3[4] DEC_X1_3[5] DEC_X1_3[6] 
+ DEC_X1_3[7] NET0133[0] NET0133[1] NET0133[2] NET0133[3] NET0133[4] 
+ NET0133[5] NET0133[6] NET0133[7] DEC_X2_3[0] DEC_X2_3[1] DEC_X2_3[2] 
+ DEC_X2_3[3] DEC_X2_3[4] DEC_X2_3[5] DEC_X2_3[6] DEC_X2_3[7] DEC_X2_SHARE_3 
+ NET0128 NET0130[0] NET0130[1] NET0130[2] NET0130[3] NET0130[4] NET0130[5] 
+ NET0130[6] NET0130[7] PD_BUF_3 NET0142 VDDHD VDDI VSSI WL_LU1[0] WL_LU1[1] 
+ WL_RU1[0] WL_RU1[1] S1AHSF400W40_SB_WLDV_U_SIM
XBK_WLDV_LD_U DEC_X0_2[0] DEC_X0_2[1] DEC_X0_2[2] DEC_X0_2[3] DEC_X0_2[4] 
+ DEC_X0_2[5] DEC_X0_2[6] DEC_X0_2[7] DEC_X0_3[0] DEC_X0_3[1] DEC_X0_3[2] 
+ DEC_X0_3[3] DEC_X0_3[4] DEC_X0_3[5] DEC_X0_3[6] DEC_X0_3[7] DEC_X1_2[0] 
+ DEC_X1_2[1] DEC_X1_2[2] DEC_X1_2[3] DEC_X1_2[4] DEC_X1_2[5] DEC_X1_2[6] 
+ DEC_X1_2[7] DEC_X1_3[0] DEC_X1_3[1] DEC_X1_3[2] DEC_X1_3[3] DEC_X1_3[4] 
+ DEC_X1_3[5] DEC_X1_3[6] DEC_X1_3[7] DEC_X2_2[0] DEC_X2_2[1] DEC_X2_2[2] 
+ DEC_X2_2[3] DEC_X2_2[4] DEC_X2_2[5] DEC_X2_2[6] DEC_X2_2[7] DEC_X2_SHARE_2 
+ DEC_X2_SHARE_3 DEC_X2_3[0] DEC_X2_3[1] DEC_X2_3[2] DEC_X2_3[3] DEC_X2_3[4] 
+ DEC_X2_3[5] DEC_X2_3[6] DEC_X2_3[7] PD_BUF_2 PD_BUF_3 VDDHD VDDI VSSI 
+ S1AHSF400W40_SB_BK_LD_U_SIM
XARR_MCB_RDR NET151 NET152 NET153 NET150 VDDI VDDHD VDDI VSSI WL_RD3[0] 
+ WL_RD3[1] WL_RD4[0] WL_RD4[1] S1AHSF400W40_SB_ARR_MCB_SIM
XARR_MCB_LUR BLB_LR_3 NET0168 BL_LR_3 NET0166 VDDI VDDHD VDDI VSSI WL_LU2[0] 
+ WL_LU2[1] WL_LU1[0] WL_LU1[1] S1AHSF400W40_SB_ARR_MCB_SIM
XARR_MCB_RUL NET171 NET516 NET173 NET170 VDDI VDDHD VDDI VSSI WL_RU1[0] 
+ WL_RU1[1] WL_RU2[0] WL_RU2[1] S1AHSF400W40_SB_ARR_MCB_SIM
XARR_MCB_RUR NET181 NET182 NET183 NET180 VDDI VDDHD VDDI VSSI WL_RU3[0] 
+ WL_RU3[1] WL_RU4[0] WL_RU4[1] S1AHSF400W40_SB_ARR_MCB_SIM
XARR_MCB_RDL NET559 NET525 NET524 NET528 VDDI VDDHD VDDI VSSI WL_RD1[0] 
+ WL_RD1[1] WL_RD2[0] WL_RD2[1] S1AHSF400W40_SB_ARR_MCB_SIM
XARR_MCB_LDL BLB_LL_1[0] BLB_LL_2 BL_LL_1[0] BL_LL_2 VDDI VDDHD VDDI VSSI 
+ WL_LD4[0] WL_LD4[1] WL_LD3[0] WL_LD3[1] S1AHSF400W40_SB_ARR_MCB_SIM
XARR_MCB_LUL BLB_LL_3 NET0218 BL_LL_3 NET0216 VDDI VDDHD VDDI VSSI WL_LU4[0] 
+ WL_LU4[1] WL_LU3[0] WL_LU3[1] S1AHSF400W40_SB_ARR_MCB_SIM
XARR_MCB_LDR BLB_LR_1[0] BLB_LR_2 BL_LR_1[0] BL_LR_2 VDDI VDDHD VDDI VSSI 
+ WL_LD2[0] WL_LD2[1] WL_LD1[0] WL_LD1[1] S1AHSF400W40_SB_ARR_MCB_SIM
XARR_BLLD_LR BLB_LR_2 BLB_LR_3 BL_LR_2 BL_LR_3 VDDI VSSI S1AHSF400W40_SB_ARR_BLLD_SIM
XARR_BLLD_LL BLB_LL_2 BLB_LL_3 BL_LL_2 BL_LL_3 VDDI VSSI S1AHSF400W40_SB_ARR_BLLD_SIM
XIO_LD_L AWT2_L3 AWT2_L2 BIST2IO_L3 BIST2IO_L2 BLEQ_L3 BLEQ_L2 CKD_L3 CKD_L2 
+ PD_BUF_L3 PD_BUF_L2 RE_L3 RE_L2 SAE_L3 SAE_L2 VDDHD VDDI VSSI WE_L3 WE_L2 
+ YL_L3[0] YL_L3[1] YL_L2[0] YL_L2[1] DEC_Y_L3[0] DEC_Y_L3[1] DEC_Y_L3[2] 
+ DEC_Y_L3[3] DEC_Y_L3[4] DEC_Y_L3[5] DEC_Y_L3[6] DEC_Y_L3[7] DEC_Y_L2[0] 
+ DEC_Y_L2[1] DEC_Y_L2[2] DEC_Y_L2[3] DEC_Y_L2[4] DEC_Y_L2[5] DEC_Y_L2[6] 
+ DEC_Y_L2[7] S1AHSF400W40_SB_IO_LD_SIM
XIO_LD_R AWT2_R2 AWT2_R3 BIST2IO_R2 BIST2IO_R3 BLEQ_R2 BLEQ_R3 CKD_R2 CKD_R3 
+ PD_BUF_R2 PD_BUF_R3 RE_R2 RE_R3 SAE_R2 SAE_R3 VDDHD VDDI VSSI WE_R2 WE_R3 
+ YL_R2[0] YL_R2[1] YL_R3[0] YL_R3[1] DEC_Y_R2[0] DEC_Y_R2[1] DEC_Y_R2[2] 
+ DEC_Y_R2[3] DEC_Y_R2[4] DEC_Y_R2[5] DEC_Y_R2[6] DEC_Y_R2[7] DEC_Y_R3[0] 
+ DEC_Y_R3[1] DEC_Y_R3[2] DEC_Y_R3[3] DEC_Y_R3[4] DEC_Y_R3[5] DEC_Y_R3[6] 
+ DEC_Y_R3[7] S1AHSF400W40_SB_IO_LD_SIM
XIO_RR AWT2_R3 AWT2_R4 BIST2IO_R3 BIST2IO_R4 NET522[0] NET522[1] NET522[2] 
+ NET522[3] NET522[4] NET522[5] NET522[6] NET522[7] NET522[8] NET522[9] 
+ NET522[10] NET522[11] NET522[12] NET522[13] NET522[14] NET522[15] NET523[0] 
+ NET523[1] NET523[2] NET523[3] NET523[4] NET523[5] NET523[6] NET523[7] 
+ NET523[8] NET523[9] NET523[10] NET523[11] NET523[12] NET523[13] NET523[14] 
+ NET523[15] BLEQ_R3 BLEQ_R4 NET519 NET520 CKD_R3 CKD_R4 NET299 NET298 
+ PD_BUF_R3 PD_BUF_R4 NET513 RE_R3 RE_R4 SAE_R3 SAE_R4 VDDHD VDDI VSSI WE_R3 
+ WE_R4 YL_R3[0] YL_R3[1] YL_R4[0] YL_R4[1] DEC_Y_R3[0] DEC_Y_R3[1] 
+ DEC_Y_R3[2] DEC_Y_R3[3] DEC_Y_R3[4] DEC_Y_R3[5] DEC_Y_R3[6] DEC_Y_R3[7] 
+ DEC_Y_R4[0] DEC_Y_R4[1] DEC_Y_R4[2] DEC_Y_R4[3] DEC_Y_R4[4] DEC_Y_R4[5] 
+ DEC_Y_R4[6] DEC_Y_R4[7] S1AHSF400W40_SB_IO_SIM
XIO_LR AWT2_L2 AWT2_L1 BIST2IO_L2 BIST2IO_L1 BL_LR_1[0] BL_LR_1[1] BL_LR_1[2] 
+ BL_LR_1[3] BL_LR_1[4] BL_LR_1[5] BL_LR_1[6] BL_LR_1[7] BL_LR_1[8] BL_LR_1[9] 
+ BL_LR_1[10] BL_LR_1[11] BL_LR_1[12] BL_LR_1[13] BL_LR_1[14] BL_LR_1[15] 
+ BLB_LR_1[0] BLB_LR_1[1] BLB_LR_1[2] BLB_LR_1[3] BLB_LR_1[4] BLB_LR_1[5] 
+ BLB_LR_1[6] BLB_LR_1[7] BLB_LR_1[8] BLB_LR_1[9] BLB_LR_1[10] BLB_LR_1[11] 
+ BLB_LR_1[12] BLB_LR_1[13] BLB_LR_1[14] BLB_LR_1[15] BLEQ_L2 BLEQ_L1 BWEB_LR 
+ BWEBM_LR CKD_L2 CKD_L1 D_LR DM_LR PD_BUF_L2 PD_BUF_L1 Q_LR RE_L2 RE_L1 
+ SAE_L2 SAE_L1 VDDHD VDDI VSSI WE_L2 WE_L1 YL_L2[0] YL_L2[1] YL_L1[0] 
+ YL_L1[1] DEC_Y_L2[0] DEC_Y_L2[1] DEC_Y_L2[2] DEC_Y_L2[3] DEC_Y_L2[4] 
+ DEC_Y_L2[5] DEC_Y_L2[6] DEC_Y_L2[7] DEC_Y_L1[0] DEC_Y_L1[1] DEC_Y_L1[2] 
+ DEC_Y_L1[3] DEC_Y_L1[4] DEC_Y_L1[5] DEC_Y_L1[6] DEC_Y_L1[7] S1AHSF400W40_SB_IO_SIM
XIO_LL AWT2_L4 AWT2_L3 BIST2IO_L4 BIST2IO_L3 BL_LL_1[0] BL_LL_1[1] BL_LL_1[2] 
+ BL_LL_1[3] BL_LL_1[4] BL_LL_1[5] BL_LL_1[6] BL_LL_1[7] BL_LL_1[8] BL_LL_1[9] 
+ BL_LL_1[10] BL_LL_1[11] BL_LL_1[12] BL_LL_1[13] BL_LL_1[14] BL_LL_1[15] 
+ BLB_LL_1[0] BLB_LL_1[1] BLB_LL_1[2] BLB_LL_1[3] BLB_LL_1[4] BLB_LL_1[5] 
+ BLB_LL_1[6] BLB_LL_1[7] BLB_LL_1[8] BLB_LL_1[9] BLB_LL_1[10] BLB_LL_1[11] 
+ BLB_LL_1[12] BLB_LL_1[13] BLB_LL_1[14] BLB_LL_1[15] BLEQ_L4 BLEQ_L3 BWEB_LL 
+ BWEBM_LL CKD_L4 CKD_L3 D_LL DM_LL PD_BUF_L4 PD_BUF_L3 Q_LL RE_L4 RE_L3 
+ SAE_L4 SAE_L3 VDDHD VDDI VSSI WE_L4 WE_L3 YL_L4[0] YL_L4[1] YL_L3[0] 
+ YL_L3[1] DEC_Y_L4[0] DEC_Y_L4[1] DEC_Y_L4[2] DEC_Y_L4[3] DEC_Y_L4[4] 
+ DEC_Y_L4[5] DEC_Y_L4[6] DEC_Y_L4[7] DEC_Y_L3[0] DEC_Y_L3[1] DEC_Y_L3[2] 
+ DEC_Y_L3[3] DEC_Y_L3[4] DEC_Y_L3[5] DEC_Y_L3[6] DEC_Y_L3[7] S1AHSF400W40_SB_IO_SIM
XIO_RL AWT2_L1 AWT2_R2 BIST2IO_L1 BIST2IO_R2 NET542[0] NET542[1] NET542[2] 
+ NET542[3] NET542[4] NET542[5] NET542[6] NET542[7] NET542[8] NET542[9] 
+ NET542[10] NET542[11] NET542[12] NET542[13] NET542[14] NET542[15] NET552[0] 
+ NET552[1] NET552[2] NET552[3] NET552[4] NET552[5] NET552[6] NET552[7] 
+ NET552[8] NET552[9] NET552[10] NET552[11] NET552[12] NET552[13] NET552[14] 
+ NET552[15] BLEQ_L1 BLEQ_R2 NET529 NET538 CKD_L1 CKD_R2 NET401 NET540 
+ PD_BUF_L1 PD_BUF_R2 NET512 RE_L1 RE_R2 SAE_L1 SAE_R2 VDDHD VDDI VSSI WE_L1 
+ WE_R2 YL_L1[0] YL_L1[1] YL_R2[0] YL_R2[1] DEC_Y_L1[0] DEC_Y_L1[1] 
+ DEC_Y_L1[2] DEC_Y_L1[3] DEC_Y_L1[4] DEC_Y_L1[5] DEC_Y_L1[6] DEC_Y_L1[7] 
+ DEC_Y_R2[0] DEC_Y_R2[1] DEC_Y_R2[2] DEC_Y_R2[3] DEC_Y_R2[4] DEC_Y_R2[5] 
+ DEC_Y_R2[6] DEC_Y_R2[7] S1AHSF400W40_SB_IO_SIM
XCNT AWT AWT2_L1 BIST BIST2IO_L1 BLEQ_L1 WL_TK CEB CEBM CKD_L1 CLK DEC_X0_1[0] 
+ DEC_X0_1[1] DEC_X0_1[2] DEC_X0_1[3] DEC_X0_1[4] DEC_X0_1[5] DEC_X0_1[6] 
+ DEC_X0_1[7] DEC_X1_1[0] DEC_X1_1[1] DEC_X1_1[2] DEC_X1_1[3] DEC_X1_1[4] 
+ DEC_X1_1[5] DEC_X1_1[6] DEC_X1_1[7] DEC_X2_1[0] DEC_X2_1[1] DEC_X2_1[2] 
+ DEC_X2_1[3] DEC_X2_1[4] DEC_X2_1[5] DEC_X2_1[6] DEC_X2_1[7] DEC_Y_L1[0] 
+ DEC_Y_L1[1] DEC_Y_L1[2] DEC_Y_L1[3] DEC_Y_L1[4] DEC_Y_L1[5] DEC_Y_L1[6] 
+ DEC_Y_L1[7] PD PD_BUF_L1 PTSEL RE_L1 RTSEL[0] RTSEL[1] SAE_L1 TK TM TRKBL 
+ VDDHD VDDI NET452 NET451 VSSI WE_L1 WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] X[0] 
+ X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL_L1[0] YL_L1[1] YM[0] YM[1] YM[2] 
+ YM[3] S1AHSF400W40_SB_CNT_SIM
XTKWL_LD VDDI TK_R2 TK_R3 VSSI WL_DUM_R2 WL_DUM_R3 WL_TK_R2 WL_TK_R3 
+ S1AHSF400W40_TKWL_LD_SIM
XTKWL_L VDDI TK TK_R2 VSSI WL_DUM_LT WL_DUM_R2 WL_TK WL_TK_R2 S1AHSF400W40_TKWL_SIM
XTKWL_R VDDI TK_R3 NET487 VSSI WL_DUM_R3 NET532 WL_TK_R3 WL_TK_LD S1AHSF400W40_TKWL_SIM
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    RESETD_F
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_RESETD_F BLTRKWLDRV CK2 CKP CKPD CKPDCLK IOSAEB RSTCK TK TRKBL VDDHD 
+ VSSI WEBXL WLP_SAE WLP_SAE_TK PTSEL RV[0] RV[1] WV[0] WV[1] WV[2]
*.PININFO CK2:I CKP:I WEBXL:I PTSEL:I RV[0]:I RV[1]:I WV[0]:I WV[1]:I WV[2]:I 
*.PININFO BLTRKWLDRV:O CKPD:O CKPDCLK:O IOSAEB:O RSTCK:O WLP_SAE:O TK:B 
*.PININFO TRKBL:B VDDHD:B VSSI:B WLP_SAE_TK:B
XTSEL_READ CKP RV[0] RV[1] VDDHD VSSI RTD_01_11 RTD_10 S1AHSF400W40_RESETD_TSEL
MP16 WLP_SAE TRKBL2 VDDHD VDDHD PCH L=60N W=2U M=4
MN7 WLP_SAE TRKBL2 VSSI VSSI NCH L=60N W=1U M=4
XI584 CKP RTD_01_11 RTD_10 VSSI VDDHD RTKB S1AHSF400W40_ANAND3 FN3=1 WN3=2U LN3=60N FN2=1 
+ WN2=2U LN2=60N FN1=1 WN1=2U LN1=60N FP1=1 WP1=1.5U LP1=60N FP2=1 WP2=1.5U 
+ LP2=60N FP3=1 WP3=1.5U LP3=60N M=1
XNAND4 TRKBL1B CKP VSSI VDDHD RSTCKB S1AHSF400W40_ANAND FN2=1 WN2=0.8U LN2=0.06U FN1=1 
+ WN1=0.8U LN1=0.06U FP1=1 WP1=0.6U LP1=0.06U FP2=1 WP2=0.6U LP2=0.06U M=1
XI592 Z6 Z5 VSSI VDDHD Z7 S1AHSF400W40_ANAND FN2=1 WN2=0.25U LN2=0.06U FN1=1 WN1=0.25U 
+ LN1=0.06U FP1=1 WP1=0.3U LP1=0.06U FP2=1 WP2=0.3U LP2=0.06U M=1
XI521 WLP_SAE3B WLP_SAE_TK1B VSSI VDDHD NET342 S1AHSF400W40_ANAND FN2=1 WN2=0.25U 
+ LN2=0.06U FN1=1 WN1=0.25U LN1=0.06U FP1=1 WP1=0.3U LP1=0.06U FP2=1 WP2=0.3U 
+ LP2=0.06U M=1
XI575 WEBXL TRKBL1B VSSI VDDHD TRKBL2 S1AHSF400W40_ANAND FN2=1 WN2=1U LN2=60N FN1=1 
+ WN1=1U LN1=60N FP1=1 WP1=1U LP1=60N FP2=1 WP2=1U LP2=60N M=2
XI589 Z3 VSSI VDDHD Z4 S1AHSF400W40_AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=0.4U LP=0.06U M=1
XI598 WLP_SAE VSSI VDDHD WLP_SAE_1B S1AHSF400W40_AINV FN=1 WN=0.4U LN=0.06U FP=1 WP=0.4U 
+ LP=0.06U M=1
XI601 WLP_SAE2 VSSI VDDHD WLP_SAE3B S1AHSF400W40_AINV FN=1 WN=0.4U LN=0.06U FP=1 WP=0.4U 
+ LP=0.06U M=1
XI620 RSTCKB VSSI VDDHD RSTCK S1AHSF400W40_AINV FN=1 WN=0.4U LN=60N FP=1 WP=0.6U LP=60N 
+ M=2
XI618 NET327 VSSI VDDHD NET299 S1AHSF400W40_AINV FN=2 WN=0.75U LN=60N FP=2 WP=1.5U LP=60N 
+ M=1
*XI585 Z0 VSSI VDDHD Z1 AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=0.4U LP=0.06U M=1
XI586 Z6 VSSI VDDHD Z0 S1AHSF400W40_AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=0.4U LP=0.06U M=1
XI606 CKPD VSSI VDDHD Z10 S1AHSF400W40_AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=0.4U LP=0.06U 
+ M=1
XI607 Z10 VSSI VDDHD CKPDCLK S1AHSF400W40_AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=0.4U 
+ LP=0.06U M=1
XI594 Z8 VSSI VDDHD CKPD S1AHSF400W40_AINV FN=8 WN=0.3U LN=0.06U FP=8 WP=0.6U LP=0.06U M=1
XI593 Z7 VSSI VDDHD Z8 S1AHSF400W40_AINV FN=2 WN=0.3U LN=0.06U FP=2 WP=0.6U LP=0.06U M=1
XI566 WLP_SAE_TK VSSI VDDHD WLP_SAE_TK1B S1AHSF400W40_AINV FN=1 WN=0.4U LN=0.06U FP=1 
+ WP=0.4U LP=0.06U M=1
XI600 WLP_SAE_1B VSSI VDDHD WLP_SAE2 S1AHSF400W40_AINV FN=1 WN=0.4U LN=0.06U FP=1 WP=0.4U 
+ LP=0.06U M=1
XI591 CKP VSSI VDDHD Z6 S1AHSF400W40_AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=0.4U LP=0.06U M=1
XI619 NET342 VSSI VDDHD NET327 S1AHSF400W40_AINV FN=1 WN=0.4U LN=60N FP=1 WP=0.8U LP=60N 
+ M=1
XI617 NET299 VSSI VDDHD IOSAEB S1AHSF400W40_AINV FN=8 WN=0.75U LN=60N FP=8 WP=1.5U LP=60N 
+ M=1
XI537 RTKB VSSI VDDHD BLTRKWLDRV S1AHSF400W40_AINV FN=6 WN=0.5U LN=60N FP=6 WP=1U LP=60N 
+ M=1
XI588 Z0 VSSI VDDHD Z3 S1AHSF400W40_AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=0.4U LP=0.06U M=1
XI590 Z4 VSSI VDDHD Z5 S1AHSF400W40_AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=0.4U LP=0.06U M=1
XI574 TRKBL VSSI VDDHD TRKBL1B S1AHSF400W40_AINV FN=1 WN=0.4U LN=60N FP=1 WP=0.8U LP=60N 
+ M=1
*XI587 Z1 VSSI VDDHD Z2 AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=0.4U LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    DECB1
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_DECB1 CKP CLK DEC EN ENC PREDEC VDDHD VSSI
*.PININFO CKP:I CLK:I EN:I ENC:I PREDEC:I DEC:O VDDHD:B VSSI:B
MM4 VDDHD PREDEC NT1 VDDHD PCH L=60N W=1.5U M=1
MM2 NET65 CKP NT1 VDDHD PCH L=60N W=1.5U M=1
MM1 VDDHD CLK NET65 VDDHD PCH L=60N W=1.5U M=1
MP0 DEC NT1 VDDHD VDDHD PCH L=60N W=2U M=6
MP5 VDDHD EN NT1 VDDHD PCH L=60N W=1.5U M=2
MN0 DEC NT1 VSSI VSSI NCH L=60N W=1U M=6
MM5 NT3 PREDEC ENC VSSI NCH L=60N W=1.5U M=2
MM0 NT1 CLK NT3 VSSI NCH L=60N W=1.5U M=2
MTN1 NT1 CKP NT3 VSSI NCH L=60N W=1.5U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    WEBBUF
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_WEBBUF BIST1B BIST2 CKC CKT VDDHD VSSI WEB WEBM WEBXL WEBXL1B
*.PININFO BIST1B:I BIST2:I CKC:I CKT:I WEB:I WEBM:I WEBXL:O WEBXL1B:O VDDHD:B 
*.PININFO VSSI:B
MM20 WEBXL CKC NET0115 VDDHD PCH L=60N W=300N M=1
MM21 NET0115 WEBXL1B VDDHD VDDHD PCH L=60N W=300N M=1
MM16 N5 CKT VDDHD VDDHD PCH L=60N W=1U M=2
MM6 WEBXL WEBX N5 VDDHD PCH L=60N W=1U M=2
MM10 WEBX WEB VDDHD VDDHD PCH L=60N W=600N M=1
MM0 WEBXL WEBX N7 VSSI NCH L=60N W=500N M=2
MM19 WEBXL CKT NET076 VSSI NCH L=60N W=300N M=1
MM18 NET076 WEBXL1B VSSI VSSI NCH L=60N W=300N M=1
MM12 WEBX WEB VSSI VSSI NCH L=60N W=300N M=1
MM17 N7 CKC VSSI VSSI NCH L=60N W=500N M=2
XI25 WEBXL VSSI VDDHD WEBXL1B S1AHSF400W40_AINV FN=2 WN=0.5U LN=0.06U FP=2 WP=1U LP=0.06U 
+ M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    AWTD
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_AWTD AWT AWT2 PD VDDHD VDDI VSSI
*.PININFO AWT:I PD:I AWT2:O VDDHD:B VDDI:B VSSI:B
XINV0 AWT1B VSSI VDDHD AWT2 S1AHSF400W40_AINV FN=12 WN=0.5U LN=0.06U FP=12 WP=1U LP=0.06U 
+ M=1
XINV1 AWT VSSI VDDHD AWT1B S1AHSF400W40_AINV FN=3 WN=0.5U LN=0.06U FP=3 WP=1U LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    BISTD
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BISTD BIST BIST1B BIST2 BIST2IO VDDHD VSSI
*.PININFO BIST:I BIST1B:O BIST2:O BIST2IO:O VDDHD:B VSSI:B
XINV2 BIST1B_2 VSSI VDDHD BIST2 S1AHSF400W40_AINV FN=3 WN=0.95U LN=0.06U FP=3 WP=1.9U 
+ LP=0.06U M=1
XINV1 BIST VSSI VDDHD BIST1B_2 S1AHSF400W40_AINV FN=1 WN=0.95U LN=0.06U FP=1 WP=1.9U 
+ LP=0.06U M=1
XINV3 BIST1B_2 VSSI VDDHD BIST2IO S1AHSF400W40_AINV FN=6 WN=0.95U LN=0.06U FP=6 WP=1.9U 
+ LP=0.06U M=1
XI21 BIST VSSI VDDHD BIST1B S1AHSF400W40_AINV FN=3 WN=0.95U LN=0.06U FP=3 WP=1.9U 
+ LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CKG
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CKG CKP CLK EN RSC RSTCK TM VDDHD VSSI
*.PININFO CLK:I EN:I RSTCK:I TM:I CKP:O RSC:O VDDHD:B VSSI:B
XINV0 Z17 VSSI VDDHD RSC S1AHSF400W40_AINV FN=2 WN=0.3U LN=0.06U FP=2 WP=0.6U LP=0.06U M=1
XNAND4 CKPC Z19 VSSI VDDHD CKP S1AHSF400W40_ANAND FN2=2 WN2=1.5U LN2=0.06U FN1=2 WN1=1.5U 
+ LN1=0.06U FP1=4 WP1=1U LP1=0.06U FP2=2 WP2=1U LP2=0.06U M=1
XNAND5 CKP RSC VSSI VDDHD Z19 S1AHSF400W40_ANAND FN2=1 WN2=0.54U LN2=0.06U FN1=1 
+ WN1=0.54U LN1=0.06U FP1=1 WP1=0.75U LP1=0.06U FP2=1 WP2=0.75U LP2=0.06U M=1
XNAND3 Z16 Z14 VSSI VDDHD Z17 S1AHSF400W40_ANAND FN2=1 WN2=0.54U LN2=0.06U FN1=1 
+ WN1=0.54U LN1=0.06U FP1=1 WP1=0.54U LP1=0.06U FP2=1 WP2=0.54U LP2=0.06U M=1
XI49 Z17 CLK VSSI VDDHD Z14 S1AHSF400W40_ANAND FN2=1 WN2=0.4U LN2=0.06U FN1=1 WN1=0.4U 
+ LN1=0.06U FP1=1 WP1=0.4U LP1=0.06U FP2=1 WP2=0.4U LP2=0.06U M=1
XI48 RSTCK Z15 VSSI VDDHD Z16 S1AHSF400W40_ANAND FN2=1 WN2=0.4U LN2=0.06U FN1=1 WN1=0.4U 
+ LN1=0.06U FP1=1 WP1=0.4U LP1=0.06U FP2=1 WP2=0.4U LP2=0.06U M=1
XNAND0 TM CLK VSSI VDDHD Z15 S1AHSF400W40_ANAND FN2=1 WN2=0.4U LN2=0.06U FN1=1 WN1=0.4U 
+ LN1=0.06U FP1=1 WP1=0.4U LP1=0.06U FP2=1 WP2=0.4U LP2=0.06U M=1
XNAND12 CLK EN RSC VSSI VDDHD CKPC S1AHSF400W40_ANAND3 FN3=1 WN3=2U LN3=0.06U FN2=1 
+ WN2=2U LN2=0.06U FN1=1 WN1=2U LN1=0.06U FP1=1 WP1=1U LP1=0.06U FP2=1 WP2=1U 
+ LP2=0.06U FP3=1 WP3=1U LP3=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    PDBUF
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_PDBUF PD PDBUF VDDI VSSI
*.PININFO PD:I PDBUF:O VDDI:B VSSI:B
XINV0 PD VSSI VDDI NET37 S1AHSF400W40_AINV FN=2 WN=0.95U LN=0.06U FP=2 WP=1.4U LP=0.06U 
+ M=1
XINV2 NET37 VSSI VDDI PDBUF S1AHSF400W40_AINV FN=8 WN=0.95U LN=0.06U FP=8 WP=1.4U 
+ LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    COTH_F
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_COTH_F AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKD CKP 
+ CKPD CLK EN ENC_D EN_D PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL 
+ VDDHD VDDI VHI VLO VSSI WEB WEBM WEBXL WEBXL1B WLP_SAE WLP_SAEB WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2]
*.PININFO AWT:I BIST:I CK1B:I CK2:I CLK:I EN:I ENC_D:I EN_D:I PD:I PTSEL:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I AWT2:O BIST1B:O BIST2:O BIST2IO:O BLTRKWLDRV:O CKD:O 
*.PININFO CKP:O CKPD:O PD_BUF:O RSC:O VHI:O VLO:O WEBXL:O WEBXL1B:O WLP_SAE:O 
*.PININFO WLP_SAEB:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE_TK:B
XRESETD BLTRKWLDRV CK2 CKP CKPD CKPDCLK WLP_SAEB RSTCK TK TRKBL VDDHD VSSI 
+ WEBXL WLP_SAE WLP_SAE_TK PTSEL RTSEL[0] RTSEL[1] WTSEL[0] WTSEL[1] WTSEL[2] 
+ S1AHSF400W40_RESETD_F
XIDEC_CKD CKPDCLK CLK CKD EN_D ENC_D WEBXL1B VDDHD VSSI S1AHSF400W40_DECB1
XWEBBUF BIST1B BIST2 CK1B CK2 VDDHD VSSI WEB WEBM WEBXL WEBXL1B S1AHSF400W40_WEBBUF
XVHILO VDDHD VHI VLO VSSI S1AHSF400W40_VHILO
XAWTD AWT AWT2 PD VDDHD VDDI VSSI S1AHSF400W40_AWTD
XBISTD BIST BIST1B BIST2 BIST2IO VDDHD VSSI S1AHSF400W40_BISTD
XCKG CKP CLK EN RSC RSTCK TM VDDHD VSSI S1AHSF400W40_CKG
XPDBUF PD PD_BUF VDDI VSSI S1AHSF400W40_PDBUF
MP2 VDDHD PD VDDI VDDI PCH L=60N W=5U M=19
MP1 VDDHD PD VDDI VDDI PCH L=60N W=3.5U M=8
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    ABUF
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ABUF A AM AX1B AX1BL AX1BL1B BIST1B BIST2 CK1B CK2 VDDHD VSSI
*.PININFO A:I AM:I BIST1B:I BIST2:I CK1B:I CK2:I AX1B:O AX1BL:O AX1BL1B:O 
*.PININFO VDDHD:B VSSI:B
MM26 AX1BL CK1B NET63 VDDHD PCH L=60N W=300N M=1
MM27 NET63 AX1BL1B VDDHD VDDHD PCH L=60N W=300N M=1
MM28 N5 CK2 VDDHD VDDHD PCH L=60N W=1U M=2
MM29 AX1BL A N5 VDDHD PCH L=60N W=1U M=2
MM19 AX1BL A N7 VSSI NCH L=60N W=500N M=2
MM20 AX1BL CK2 NET84 VSSI NCH L=60N W=300N M=1
MM21 NET84 AX1BL1B VSSI VSSI NCH L=60N W=300N M=1
MM23 N7 CK1B VSSI VSSI NCH L=60N W=500N M=2
XI25 AX1BL VSSI VDDHD AX1BL1B S1AHSF400W40_AINV FN=2 WN=0.5U LN=0.06U FP=2 WP=1U LP=0.06U 
+ M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    DECB1YL
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_DECB1YL CKP CLK DEC EN ENC PREDEC VDDHD VSSI
*.PININFO CKP:I CLK:I EN:I ENC:I PREDEC:I DEC:O VDDHD:B VSSI:B
MP0 DEC NT1 VDDHD VDDHD PCH L=60N W=2U M=9
MM3 VDDHD PREDEC NT1 VDDHD PCH L=60N W=1.2U M=1
MN0 DEC NT1 VSSI VSSI NCH L=60N W=1U M=9
MTN2 NT1 PREDEC VSSI VSSI NCH L=60N W=1.4U M=5
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    DECB4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_DECB4 IN0A IN0B IN1A IN1B IN2 PREDEC0 PREDEC1 PREDEC2 PREDEC3 VDDHD 
+ VSSI
*.PININFO IN0A:I IN0B:I IN1A:I IN1B:I IN2:I PREDEC0:O PREDEC1:O PREDEC2:O 
*.PININFO PREDEC3:O VDDHD:B VSSI:B
MM1 NET0134 IN0A VDDHD VDDHD PCH L=60N W=400N M=1
MM2 NET0134 IN1A VDDHD VDDHD PCH L=60N W=400N M=1
MM4 NET0138 IN0B VDDHD VDDHD PCH L=60N W=400N M=1
MM5 NET0138 IN1A VDDHD VDDHD PCH L=60N W=400N M=1
MM25 NET0134 IN2 VDDHD VDDHD PCH L=60N W=400N M=2
MM24 NET0138 IN2 VDDHD VDDHD PCH L=60N W=400N M=2
MM23 NET0154 IN2 VDDHD VDDHD PCH L=60N W=400N M=2
MM22 NET0150 IN2 VDDHD VDDHD PCH L=60N W=400N M=2
MM18 NET0150 IN0A VDDHD VDDHD PCH L=60N W=400N M=1
MM17 NET0150 IN1B VDDHD VDDHD PCH L=60N W=400N M=1
MM16 NET0154 IN0B VDDHD VDDHD PCH L=60N W=400N M=1
MM15 NET0154 IN1B VDDHD VDDHD PCH L=60N W=400N M=1
MM3 N2 IN1A NET19 VSSI NCH L=60N W=600N M=1
MM6 N5 IN1B NET19 VSSI NCH L=60N W=600N M=1
MM0 NET0134 IN0A N2 VSSI NCH L=60N W=600N M=1
MM7 NET0138 IN0B NET0179 VSSI NCH L=60N W=600N M=1
MM8 NET0179 IN1A NET19 VSSI NCH L=60N W=600N M=1
MM26 NET19 IN2 VSSI VSSI NCH L=60N W=600N M=4
MM21 NET0150 IN0A N5 VSSI NCH L=60N W=600N M=1
MM20 NET0154 IN0B NET0199 VSSI NCH L=60N W=600N M=1
MM19 NET0199 IN1B NET19 VSSI NCH L=60N W=600N M=1
XINV0 NET0134 VSSI VDDHD PREDEC0 S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=0.8U 
+ LP=0.06U M=1
XINV1 NET0138 VSSI VDDHD PREDEC1 S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=0.8U 
+ LP=0.06U M=1
XINV2 NET0150 VSSI VDDHD PREDEC2 S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=0.8U 
+ LP=0.06U M=1
XINV3 NET0154 VSSI VDDHD PREDEC3 S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=0.8U 
+ LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    DECB2
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_DECB2 IN0A IN0B IN1 PREDEC0 PREDEC1 VDDHD VSSI
*.PININFO IN0A:I IN0B:I IN1:I PREDEC0:O PREDEC1:O VDDHD:B VSSI:B
MM4 N3 IN0B VDDHD VDDHD PCH L=60N W=400N M=1
MM5 N3 IN1 VDDHD VDDHD PCH L=60N W=400N M=2
MM1 N1 IN0A VDDHD VDDHD PCH L=60N W=400N M=1
MM2 N1 IN1 VDDHD VDDHD PCH L=60N W=400N M=2
MM3 NET70 IN1 VSSI VSSI NCH L=60N W=600N M=1
MM8 NET75 IN1 VSSI VSSI NCH L=60N W=600N M=1
MM7 N3 IN0B NET75 VSSI NCH L=60N W=600N M=1
MM0 N1 IN0A NET70 VSSI NCH L=60N W=600N M=1
XINV1 N1 VSSI VDDHD PREDEC0 S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U LP=0.06U 
+ M=1
XINV0 N3 VSSI VDDHD PREDEC1 S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U LP=0.06U 
+ M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CKBUF
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CKBUF CK1B CK2 CKP CLK VDDHD VSSI
*.PININFO CKP:I CLK:I CK1B:O CK2:O VDDHD:B VSSI:B
XINV0 CK1B VSSI VDDHD CK2 S1AHSF400W40_AINV FN=6 WN=0.75U LN=0.06U FP=6 WP=1.5U LP=0.06U 
+ M=1
XNOR0 CKP CLK VSSI VDDHD CK1B S1AHSF400W40_ANOR FN2=4 WN2=0.9U LN2=0.06U FN1=1 WN1=0.5U 
+ LN1=0.06U FP1=3 WP1=1.5U LP1=0.06U FP2=3 WP2=1.5U LP2=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    ENBUFB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ENBUFB BIST1B BIST2 CEB CEBM CK1B CK2 EN ENC ENC_XY ENC_Z EN_D EN_DCLK 
+ RSC VDDHD VSSI
*.PININFO BIST1B:I BIST2:I CEB:I CEBM:I CK1B:I CK2:I RSC:I EN:O ENC:O ENC_XY:O 
*.PININFO ENC_Z:O EN_D:O EN_DCLK:O VDDHD:B VSSI:B
MM1 CEBXL CK1B NET0203 VDDHD PCH L=60N W=500N M=1
MM16 CEBXL CEBX N5 VDDHD PCH L=60N W=1U M=2
MM7 CEBXL RSC VDDHD VDDHD PCH L=60N W=1.4U M=1
MM2 NET0203 EN VDDHD VDDHD PCH L=60N W=500N M=1
MM19 N5 CK2 VDDHD VDDHD PCH L=60N W=1U M=2
MM10 CEBX CEB VDDHD VDDHD PCH L=60N W=500N M=1
MN300 ENC EN VSSI VSSI NCH L=60N W=2U M=4
MM18 N7 CK1B NET0151 VSSI NCH L=60N W=1U M=1
MM17 CEBXL CEBX N7 VSSI NCH L=60N W=1U M=1
MM20 NET0151 RSC VSSI VSSI NCH L=60N W=1U M=2
MM3 CEBXL CK2 NET0168 VSSI NCH L=60N W=500N M=1
MM4 NET0168 EN NET0188 VSSI NCH L=60N W=500N M=1
MN200 ENC_Z EN VSSI VSSI NCH L=60N W=2U M=4
MM5 NET0188 RSC VSSI VSSI NCH L=60N W=1U M=1
MN100 ENC_XY EN VSSI VSSI NCH L=60N W=2U M=4
MM12 CEBX CEB VSSI VSSI NCH L=60N W=500N M=1
XI141 CEBXL VSSI VDDHD EN S1AHSF400W40_AINV FN=2 WN=2U LN=0.06U FP=6 WP=1.4U LP=0.06U M=1
XI161 NET122 VSSI VDDHD EN_DCLK S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U 
+ LP=0.06U M=1
XI162 NET100 VSSI VDDHD NET0240 S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U 
+ LP=0.06U M=1
XINV5 NET0240 VSSI VDDHD NET94 S1AHSF400W40_AINV FN=3 WN=0.5U LN=0.06U FP=3 WP=1U 
+ LP=0.06U M=1
XI152 NET94 VSSI VDDHD EN_D S1AHSF400W40_AINV FN=6 WN=0.75U LN=0.06U FP=6 WP=1.6U 
+ LP=0.06U M=1
XINV10 NET112 VSSI VDDHD NET103 S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.3U 
+ LP=0.06U M=1
XINV8 NET115 VSSI VDDHD NET109 S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.3U 
+ LP=0.06U M=1
XINV9 NET109 VSSI VDDHD NET112 S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.3U 
+ LP=0.06U M=1
XINV7 EN VSSI VDDHD NET115 S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.3U LP=0.06U 
+ M=1
XI158 NET103 EN VSSI VDDHD NET100 S1AHSF400W40_ANOR FN2=1 WN2=0.3U LN2=0.06U FN1=1 
+ WN1=0.3U LN1=0.06U FP1=1 WP1=0.6U LP1=0.06U FP2=1 WP2=0.6U LP2=0.06U M=1
XNOR0 EN EN VSSI VDDHD NET122 S1AHSF400W40_ANOR FN2=1 WN2=0.3U LN2=0.06U FN1=1 WN1=0.3U 
+ LN1=0.06U FP1=1 WP1=0.6U LP1=0.06U FP2=1 WP2=0.6U LP2=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CDEC_M8M16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CDEC_M8M16 AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8] AX[9] 
+ AX[10] BIST1B BIST2 CEB CEBM CK1B CK2 CKP CKPD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] 
+ DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN ENC EN_DCLK PD REDEN REDENB 
+ RSC RW_RE VDDHD VDDI VSSI WEBXL WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] 
+ X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] 
+ XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO BIST1B:I BIST2:I CEB:I CEBM:I CKP:I CKPD:I CLK:I PD:I REDEN:I 
*.PININFO REDENB:I RSC:I WEBXL:I WEBXL1B:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I 
*.PININFO X[5]:I X[6]:I X[7]:I X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I 
*.PININFO XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I 
*.PININFO Y[0]:I Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AX[0]:O 
*.PININFO AX[1]:O AX[2]:O AX[3]:O AX[4]:O AX[5]:O AX[6]:O AX[7]:O AX[8]:O 
*.PININFO AX[9]:O AX[10]:O CK1B:O CK2:O DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O 
*.PININFO DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O 
*.PININFO DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O 
*.PININFO DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O 
*.PININFO DEC_X2[2]:O DEC_X2[3]:O DEC_X3[0]:O DEC_X3[1]:O DEC_X3[2]:O 
*.PININFO DEC_X3[3]:O DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O DEC_X3[7]:O 
*.PININFO DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O DEC_Y[5]:O 
*.PININFO DEC_Y[6]:O DEC_Y[7]:O EN:O ENC:O EN_DCLK:O RW_RE:O YL[0]:O VDDHD:B 
*.PININFO VDDI:B VSSI:B
XABUF_Y<2> Y[2] YM[2] NET140 AYC[2] AYT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_X<3> X[3] XM[3] AX[3] AXC[3] AXT[3] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_X<4> X[4] XM[4] AX[4] AXC[4] AXT[4] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_X<5> X[5] XM[5] AX[5] AXC[5] AXT[5] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_X<8> X[8] XM[8] AX[8] AXC[8] AXT[8] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_X<9> X[9] XM[9] AX[9] AXC[9] AXT[9] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_X<10> X[10] XM[10] AX[10] AXC[10] AXT[10] BIST1B BIST2 CK1B CK2 VDDHD 
+ VSSI S1AHSF400W40_ABUF
XABUF_X<0> X[0] XM[0] AX[0] AXC[0] AXT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_X<1> X[1] XM[1] AX[1] AXC[1] AXT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_X<2> X[2] XM[2] AX[2] AXC[2] AXT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_Y<0> Y[0] YM[0] NET123[0] AYC[0] AYT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_Y<1> Y[1] YM[1] NET123[1] AYC[1] AYT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_X<6> X[6] XM[6] AX[6] AXC[6] AXT[6] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_X<7> X[7] XM[7] AX[7] AXC[7] AXT[7] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_Y<3> Y[3] YM[3] NET206 NET204 AYT[3] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XIDEC_YL CKPD CLK YL[0] EN_D ENC_XY AYT[3] VDDHD VSSI S1AHSF400W40_DECB1YL
XIPDEC_X0<0> AXC[0] AXT[0] AXC[1] AXT[1] AXC[2] XA[0] XA[1] XA[2] XA[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_X0<1> AXC[0] AXT[0] AXC[1] AXT[1] AXT[2] XA[4] XA[5] XA[6] XA[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_X3<0> AXC[8] AXT[8] AXC[9] AXT[9] AXC[10] Z[0] Z[1] Z[2] Z[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_X3<1> AXC[8] AXT[8] AXC[9] AXT[9] AXT[10] Z[4] Z[5] Z[6] Z[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_X1<0> AXC[3] AXT[3] AXC[4] AXT[4] AXC[5] XB[0] XB[1] XB[2] XB[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_X1<1> AXC[3] AXT[3] AXC[4] AXT[4] AXT[5] XB[4] XB[5] XB[6] XB[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_Y<0> AYC[0] AYT[0] AYC[1] AYT[1] AYC[2] XY[0] XY[1] XY[2] XY[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_Y<1> AYC[0] AYT[0] AYC[1] AYT[1] AYT[2] XY[4] XY[5] XY[6] XY[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIDEC_X0<0> CKPD CLK DEC_X0[0] EN_D ENC XA[0] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<1> CKPD CLK DEC_X0[1] EN_D ENC XA[1] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<2> CKPD CLK DEC_X0[2] EN_D ENC XA[2] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<3> CKPD CLK DEC_X0[3] EN_D ENC XA[3] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<4> CKPD CLK DEC_X0[4] EN_D ENC XA[4] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<5> CKPD CLK DEC_X0[5] EN_D ENC XA[5] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<6> CKPD CLK DEC_X0[6] EN_D ENC XA[6] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<7> CKPD CLK DEC_X0[7] EN_D ENC XA[7] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_RWRE CKPD CLK RW_RE EN_D ENC_XY WEBXL VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<0> CKPD CLK DEC_Y[0] EN_D ENC_XY XY[0] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<1> CKPD CLK DEC_Y[1] EN_D ENC_XY XY[1] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<2> CKPD CLK DEC_Y[2] EN_D ENC_XY XY[2] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<3> CKPD CLK DEC_Y[3] EN_D ENC_XY XY[3] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<0> CKP CLK DEC_X3[0] EN ENC_Z Z[0] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<1> CKP CLK DEC_X3[1] EN ENC_Z Z[1] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<2> CKP CLK DEC_X3[2] EN ENC_Z Z[2] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<3> CKP CLK DEC_X3[3] EN ENC_Z Z[3] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<4> CKP CLK DEC_X3[4] EN ENC_Z Z[4] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<5> CKP CLK DEC_X3[5] EN ENC_Z Z[5] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<6> CKP CLK DEC_X3[6] EN ENC_Z Z[6] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<7> CKP CLK DEC_X3[7] EN ENC_Z Z[7] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<4> CKPD CLK DEC_Y[4] EN_D ENC_XY XY[4] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<5> CKPD CLK DEC_Y[5] EN_D ENC_XY XY[5] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<6> CKPD CLK DEC_Y[6] EN_D ENC_XY XY[6] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<7> CKPD CLK DEC_Y[7] EN_D ENC_XY XY[7] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X2<0> CKPD CLK DEC_X2[0] EN_D ENC_XY XC[0] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X2<1> CKPD CLK DEC_X2[1] EN_D ENC_XY XC[1] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X2<2> CKPD CLK DEC_X2[2] EN_D ENC_XY XC[2] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X2<3> CKPD CLK DEC_X2[3] EN_D ENC_XY XC[3] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<0> CKPD CLK DEC_X1[0] EN_D ENC XB[0] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<1> CKPD CLK DEC_X1[1] EN_D ENC XB[1] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<2> CKPD CLK DEC_X1[2] EN_D ENC XB[2] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<3> CKPD CLK DEC_X1[3] EN_D ENC XB[3] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<4> CKPD CLK DEC_X1[4] EN_D ENC XB[4] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<5> CKPD CLK DEC_X1[5] EN_D ENC XB[5] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<6> CKPD CLK DEC_X1[6] EN_D ENC XB[6] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<7> CKPD CLK DEC_X1[7] EN_D ENC XB[7] VDDHD VSSI S1AHSF400W40_DECB1
XIPDEC_X2<0> AXC[6] AXT[6] AXC[7] XC[0] XC[1] VDDHD VSSI S1AHSF400W40_DECB2
XIPDEC_X2<1> AXC[6] AXT[6] AXT[7] XC[2] XC[3] VDDHD VSSI S1AHSF400W40_DECB2
XCKBUF CK1B CK2 CKPD CLK VDDHD VSSI S1AHSF400W40_CKBUF
XCEBBUF BIST1B BIST2 CEB CEBM CK1B CK2 EN ENC ENC_XY ENC_Z EN_D EN_DCLK RSC 
+ VDDHD VSSI S1AHSF400W40_ENBUFB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_F_M16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_F_M16 AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD 
+ PD_BUF PD_CVDDBUF PTSEL REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL 
+ VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] 
+ WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] 
+ XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] 
+ Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I REDEN:I REDENB:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I 
*.PININFO XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I 
*.PININFO Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O BIST2IO:O 
*.PININFO BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O 
*.PININFO DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O DEC_X1[0]:O 
*.PININFO DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O DEC_X1[5]:O 
*.PININFO DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O DEC_X2[2]:O 
*.PININFO DEC_X2[3]:O DEC_X3[0]:O DEC_X3[1]:O DEC_X3[2]:O DEC_X3[3]:O 
*.PININFO DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O DEC_X3[7]:O DEC_Y[0]:O 
*.PININFO DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O 
*.PININFO DEC_Y[7]:O PD_BUF:O PD_CVDDBUF:O RW_RE:O VHI:O VLO:O WLP_SAE:O 
*.PININFO WLP_SAEB:O YL[0]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE_TK:B
XCOTHERS AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKD CKP CKPD 
+ CLK EN ENC EN_DCLK PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WEB WEBM WEBXL WEBXL1B WLP_SAE WLP_SAEB WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2] S1AHSF400W40_COTH_F
XCDEC AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8] AX[9] AX[10] 
+ BIST1B BIST2 CEB CEBM CK1B CK2 CKP CKPD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN ENC EN_DCLK PD REDEN REDENB RSC RW_RE 
+ VDDHD VDDI VSSI WEBXL WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] 
+ X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] 
+ XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3] S1AHSF400W40_CDEC_M8M16
MX0_PD<0> DEC_X0[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<1> DEC_X0[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<2> DEC_X0[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<3> DEC_X0[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<4> DEC_X0[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<5> DEC_X0[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<6> DEC_X0[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<7> DEC_X0[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<0> DEC_X1[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<1> DEC_X1[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<2> DEC_X1[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<3> DEC_X1[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<4> DEC_X1[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<5> DEC_X1[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<6> DEC_X1[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<7> DEC_X1[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_F_M8
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_F_M8 AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD 
+ PD_BUF PD_CVDDBUF PTSEL REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL 
+ VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] 
+ WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] 
+ XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] 
+ Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I REDEN:I REDENB:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I 
*.PININFO XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I 
*.PININFO Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O BIST2IO:O 
*.PININFO BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O 
*.PININFO DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O DEC_X1[0]:O 
*.PININFO DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O DEC_X1[5]:O 
*.PININFO DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O DEC_X2[2]:O 
*.PININFO DEC_X2[3]:O DEC_X3[0]:O DEC_X3[1]:O DEC_X3[2]:O DEC_X3[3]:O 
*.PININFO DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O DEC_X3[7]:O DEC_Y[0]:O 
*.PININFO DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O 
*.PININFO DEC_Y[7]:O PD_BUF:O PD_CVDDBUF:O RW_RE:O VHI:O VLO:O WLP_SAE:O 
*.PININFO WLP_SAEB:O YL[0]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE_TK:B
XCOTHERS AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKD CKP CKPD 
+ CLK EN ENC EN_DCLK PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WEB WEBM WEBXL WEBXL1B WLP_SAE WLP_SAEB WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2] S1AHSF400W40_COTH_F
MX0_PD<0> DEC_X0[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<1> DEC_X0[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<2> DEC_X0[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<3> DEC_X0[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<4> DEC_X0[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<5> DEC_X0[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<6> DEC_X0[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<7> DEC_X0[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<0> DEC_X1[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<1> DEC_X1[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<2> DEC_X1[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<3> DEC_X1[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<4> DEC_X1[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<5> DEC_X1[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<6> DEC_X1[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<7> DEC_X1[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
XCDEC AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8] AX[9] AX[10] 
+ BIST1B BIST2 CEB CEBM CK1B CK2 CKP CKPD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN ENC EN_DCLK PD REDEN REDENB RSC RW_RE 
+ VDDHD VDDI VSSI WEBXL WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] 
+ X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] 
+ XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3] S1AHSF400W40_CDEC_M8M16
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CDEC_M4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CDEC_M4 AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8] AX[9] 
+ AX[10] BIST1B BIST2 CEB CEBM CK1B CK2 CKP CKPD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] 
+ DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN ENC EN_DCLK PD REDEN REDENB 
+ RSC RW_RE VDDHD VDDI VSSI WEBXL WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] 
+ X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] 
+ XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO BIST1B:I BIST2:I CEB:I CEBM:I CKP:I CKPD:I CLK:I PD:I REDEN:I 
*.PININFO REDENB:I RSC:I WEBXL:I WEBXL1B:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I 
*.PININFO X[5]:I X[6]:I X[7]:I X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I 
*.PININFO XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I 
*.PININFO Y[0]:I Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AX[0]:O 
*.PININFO AX[1]:O AX[2]:O AX[3]:O AX[4]:O AX[5]:O AX[6]:O AX[7]:O AX[8]:O 
*.PININFO AX[9]:O AX[10]:O CK1B:O CK2:O DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O 
*.PININFO DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O 
*.PININFO DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O 
*.PININFO DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O 
*.PININFO DEC_X2[2]:O DEC_X2[3]:O DEC_X3[0]:O DEC_X3[1]:O DEC_X3[2]:O 
*.PININFO DEC_X3[3]:O DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O DEC_X3[7]:O 
*.PININFO DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O DEC_Y[5]:O 
*.PININFO DEC_Y[6]:O DEC_Y[7]:O EN:O ENC:O EN_DCLK:O RW_RE:O YL[0]:O VDDHD:B 
*.PININFO VDDI:B VSSI:B
XIDEC_YL CKPD CLK YL[0] EN_D ENC_XY AYT[3] VDDHD VSSI S1AHSF400W40_DECB1YL
XCEBBUF BIST1B BIST2 CEB CEBM CK1B CK2 EN ENC ENC_XY ENC_Z EN_D EN_DCLK RSC 
+ VDDHD VSSI S1AHSF400W40_ENBUFB
XCKBUF CK1B CK2 CKPD CLK VDDHD VSSI S1AHSF400W40_CKBUF
XIPDEC_X2<0> AXC[6] AXT[6] AXC[7] XC[0] XC[1] VDDHD VSSI S1AHSF400W40_DECB2
XIPDEC_X2<1> AXC[6] AXT[6] AXT[7] XC[2] XC[3] VDDHD VSSI S1AHSF400W40_DECB2
XIDEC_X3<0> CKP CLK DEC_X3[0] EN ENC_Z Z[0] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<1> CKP CLK DEC_X3[1] EN ENC_Z Z[1] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<2> CKP CLK DEC_X3[2] EN ENC_Z Z[2] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<3> CKP CLK DEC_X3[3] EN ENC_Z Z[3] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<4> CKP CLK DEC_X3[4] EN ENC_Z Z[4] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<5> CKP CLK DEC_X3[5] EN ENC_Z Z[5] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<6> CKP CLK DEC_X3[6] EN ENC_Z Z[6] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<7> CKP CLK DEC_X3[7] EN ENC_Z Z[7] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X2<0> CKPD CLK DEC_X2[0] EN_D ENC_XY XC[0] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X2<1> CKPD CLK DEC_X2[1] EN_D ENC_XY XC[1] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X2<2> CKPD CLK DEC_X2[2] EN_D ENC_XY XC[2] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X2<3> CKPD CLK DEC_X2[3] EN_D ENC_XY XC[3] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<0> CKPD CLK DEC_X1[0] EN_D ENC XB[0] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<1> CKPD CLK DEC_X1[1] EN_D ENC XB[1] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<2> CKPD CLK DEC_X1[2] EN_D ENC XB[2] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<3> CKPD CLK DEC_X1[3] EN_D ENC XB[3] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<4> CKPD CLK DEC_X1[4] EN_D ENC XB[4] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<5> CKPD CLK DEC_X1[5] EN_D ENC XB[5] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<6> CKPD CLK DEC_X1[6] EN_D ENC XB[6] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<7> CKPD CLK DEC_X1[7] EN_D ENC XB[7] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<0> CKPD CLK DEC_X0[0] EN_D ENC XA[0] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<1> CKPD CLK DEC_X0[1] EN_D ENC XA[1] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<2> CKPD CLK DEC_X0[2] EN_D ENC XA[2] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<3> CKPD CLK DEC_X0[3] EN_D ENC XA[3] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<4> CKPD CLK DEC_X0[4] EN_D ENC XA[4] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<5> CKPD CLK DEC_X0[5] EN_D ENC XA[5] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<6> CKPD CLK DEC_X0[6] EN_D ENC XA[6] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<7> CKPD CLK DEC_X0[7] EN_D ENC XA[7] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_RWRE CKPD CLK RW_RE EN_D ENC_XY WEBXL VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<4> CKPD CLK DEC_Y[4] EN_D ENC_XY XY[4] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<5> CKPD CLK DEC_Y[5] EN_D ENC_XY XY[5] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<6> CKPD CLK DEC_Y[6] EN_D ENC_XY XY[6] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<7> CKPD CLK DEC_Y[7] EN_D ENC_XY XY[7] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<0> CKPD CLK DEC_Y[0] EN_D ENC_XY XY[0] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<1> CKPD CLK DEC_Y[1] EN_D ENC_XY XY[1] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<2> CKPD CLK DEC_Y[2] EN_D ENC_XY XY[2] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<3> CKPD CLK DEC_Y[3] EN_D ENC_XY XY[3] VDDHD VSSI S1AHSF400W40_DECB1
XIPDEC_X0<0> AXC[0] AXT[0] AXC[1] AXT[1] AXC[2] XA[0] XA[1] XA[2] XA[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_X0<1> AXC[0] AXT[0] AXC[1] AXT[1] AXT[2] XA[4] XA[5] XA[6] XA[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_Y<0> AYC[0] AYT[0] AYC[1] AYT[1] WEBXL XY[0] XY[1] XY[2] XY[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_Y<1> AYC[0] AYT[0] AYC[1] AYT[1] WEBXL1B XY[4] XY[5] XY[6] XY[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_X3<0> AXC[8] AXT[8] AXC[9] AXT[9] AXC[10] Z[0] Z[1] Z[2] Z[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_X3<1> AXC[8] AXT[8] AXC[9] AXT[9] AXT[10] Z[4] Z[5] Z[6] Z[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_X1<0> AXC[3] AXT[3] AXC[4] AXT[4] AXC[5] XB[0] XB[1] XB[2] XB[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_X1<1> AXC[3] AXT[3] AXC[4] AXT[4] AXT[5] XB[4] XB[5] XB[6] XB[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XABUF_X<6> X[6] XM[6] AX[6] AXC[6] AXT[6] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_X<7> X[7] XM[7] AX[7] AXC[7] AXT[7] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_Y<3> Y[3] YM[3] NET0283 NET207 AYT[3] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_Y<2> Y[2] YM[2] NET0294 NET217 NET216 BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_X<3> X[3] XM[3] AX[3] AXC[3] AXT[3] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_X<4> X[4] XM[4] AX[4] AXC[4] AXT[4] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_X<5> X[5] XM[5] AX[5] AXC[5] AXT[5] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_X<8> X[8] XM[8] AX[8] AXC[8] AXT[8] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_X<9> X[9] XM[9] AX[9] AXC[9] AXT[9] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_X<10> X[10] XM[10] AX[10] AXC[10] AXT[10] BIST1B BIST2 CK1B CK2 VDDHD 
+ VSSI S1AHSF400W40_ABUF
XABUF_X<0> X[0] XM[0] AX[0] AXC[0] AXT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_X<1> X[1] XM[1] AX[1] AXC[1] AXT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_X<2> X[2] XM[2] AX[2] AXC[2] AXT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_Y<0> Y[0] YM[0] NET089[0] AYC[0] AYT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
XABUF_Y<1> Y[1] YM[1] NET089[1] AYC[1] AYT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_F_M4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_F_M4 AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD 
+ PD_BUF PD_CVDDBUF PTSEL REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL 
+ VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] 
+ WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] 
+ XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] 
+ Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I REDEN:I REDENB:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I 
*.PININFO XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I 
*.PININFO Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O BIST2IO:O 
*.PININFO BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O 
*.PININFO DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O DEC_X1[0]:O 
*.PININFO DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O DEC_X1[5]:O 
*.PININFO DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O DEC_X2[2]:O 
*.PININFO DEC_X2[3]:O DEC_X3[0]:O DEC_X3[1]:O DEC_X3[2]:O DEC_X3[3]:O 
*.PININFO DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O DEC_X3[7]:O DEC_Y[0]:O 
*.PININFO DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O 
*.PININFO DEC_Y[7]:O PD_BUF:O PD_CVDDBUF:O RW_RE:O VHI:O VLO:O WLP_SAE:O 
*.PININFO WLP_SAEB:O YL[0]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE_TK:B
XCOTHERS AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKD CKP CKPD 
+ CLK EN ENC EN_DCLK PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WEB WEBM WEBXL WEBXL1B WLP_SAE WLP_SAEB WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2] S1AHSF400W40_COTH_F
MX0_PD<0> DEC_X0[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<1> DEC_X0[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<2> DEC_X0[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<3> DEC_X0[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<4> DEC_X0[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<5> DEC_X0[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<6> DEC_X0[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<7> DEC_X0[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<0> DEC_X1[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<1> DEC_X1[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<2> DEC_X1[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<3> DEC_X1[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<4> DEC_X1[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<5> DEC_X1[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<6> DEC_X1[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<7> DEC_X1[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
XCDEC AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8] AX[9] AX[10] 
+ BIST1B BIST2 CEB CEBM CK1B CK2 CKP CKPD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN ENC EN_DCLK PD REDEN REDENB RSC RW_RE 
+ VDDHD VDDI VSSI WEBXL WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] 
+ X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] 
+ XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3] S1AHSF400W40_CDEC_M4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    WEBBUF_BIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_WEBBUF_BIST BIST1B BIST2 CKC CKT VDDHD VSSI WEB WEBM WEBXL WEBXL1B
*.PININFO BIST1B:I BIST2:I CKC:I CKT:I WEB:I WEBM:I WEBXL:O WEBXL1B:O VDDHD:B 
*.PININFO VSSI:B
MM14 WEBX BIST1B N3 VDDHD PCH L=60N W=600N M=1
MM15 N3 WEBM VDDHD VDDHD PCH L=60N W=600N M=1
MM20 WEBXL CKC NET0115 VDDHD PCH L=60N W=300N M=1
MM21 NET0115 WEBXL1B VDDHD VDDHD PCH L=60N W=300N M=1
MM16 N5 CKT VDDHD VDDHD PCH L=60N W=1U M=2
MM6 WEBXL WEBX N5 VDDHD PCH L=60N W=1U M=2
MM8 WEBX BIST2 N1 VDDHD PCH L=60N W=600N M=1
MM10 N1 WEB VDDHD VDDHD PCH L=60N W=600N M=1
MM9 WEBX BIST1B N2 VSSI NCH L=60N W=300N M=1
MM11 N4 WEBM VSSI VSSI NCH L=60N W=300N M=1
MM13 WEBX BIST2 N4 VSSI NCH L=60N W=300N M=1
MM0 WEBXL WEBX N7 VSSI NCH L=60N W=500N M=2
MM19 WEBXL CKT NET076 VSSI NCH L=60N W=300N M=1
MM18 NET076 WEBXL1B VSSI VSSI NCH L=60N W=300N M=1
MM12 N2 WEB VSSI VSSI NCH L=60N W=300N M=1
MM17 N7 CKC VSSI VSSI NCH L=60N W=500N M=2
XI25 WEBXL VSSI VDDHD WEBXL1B S1AHSF400W40_AINV FN=2 WN=0.5U LN=0.06U FP=2 WP=1U LP=0.06U 
+ M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    COTH_F_BIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_COTH_F_BIST AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKD 
+ CKP CKPD CLK EN ENC_D EN_D PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL 
+ VDDHD VDDI VHI VLO VSSI WEB WEBM WEBXL WEBXL1B WLP_SAE WLP_SAEB WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2]
*.PININFO AWT:I BIST:I CK1B:I CK2:I CLK:I EN:I ENC_D:I EN_D:I PD:I PTSEL:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I AWT2:O BIST1B:O BIST2:O BIST2IO:O BLTRKWLDRV:O CKD:O 
*.PININFO CKP:O CKPD:O PD_BUF:O RSC:O VHI:O VLO:O WEBXL:O WEBXL1B:O WLP_SAE:O 
*.PININFO WLP_SAEB:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE_TK:B
XRESETD BLTRKWLDRV CK2 CKP CKPD CKPDCLK WLP_SAEB RSTCK TK TRKBL VDDHD VSSI 
+ WEBXL WLP_SAE WLP_SAE_TK PTSEL RTSEL[0] RTSEL[1] WTSEL[0] WTSEL[1] WTSEL[2] 
+ S1AHSF400W40_RESETD_F
XVHILO_SB VDDHD VHI VLO VSSI S1AHSF400W40_VHILO_SB
XWEBBUF BIST1B BIST2 CK1B CK2 VDDHD VSSI WEB WEBM WEBXL WEBXL1B S1AHSF400W40_WEBBUF_BIST
XIDEC_CKD CKPDCLK CLK CKD EN_D ENC_D WEBXL1B VDDHD VSSI S1AHSF400W40_DECB1
XAWTD AWT AWT2 PD VDDHD VDDI VSSI S1AHSF400W40_AWTD
XBISTD BIST BIST1B BIST2 BIST2IO VDDHD VSSI S1AHSF400W40_BISTD
XCKG CKP CLK EN RSC RSTCK TM VDDHD VSSI S1AHSF400W40_CKG
XPDBUF PD PD_BUF VDDI VSSI S1AHSF400W40_PDBUF
MP2 VDDHD PD VDDI VDDI PCH L=60N W=5U M=19
MP1 VDDHD PD VDDI VDDI PCH L=60N W=3.5U M=8
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    ENBUFB_BIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ENBUFB_BIST BIST1B BIST2 CEB CEBM CK1B CK2 EN ENC ENC_XY ENC_Z EN_D 
+ EN_DCLK RSC VDDHD VSSI
*.PININFO BIST1B:I BIST2:I CEB:I CEBM:I CK1B:I CK2:I RSC:I EN:O ENC:O ENC_XY:O 
*.PININFO ENC_Z:O EN_D:O EN_DCLK:O VDDHD:B VSSI:B
MM1 CEBXL CK1B NET0203 VDDHD PCH L=60N W=500N M=1
MM16 CEBXL CEBX N5 VDDHD PCH L=60N W=1U M=2
MM7 CEBXL RSC VDDHD VDDHD PCH L=60N W=1.4U M=1
MM15 NET0135 CEBM VDDHD VDDHD PCH L=60N W=500N M=1
MM2 NET0203 EN VDDHD VDDHD PCH L=60N W=500N M=1
MM19 N5 CK2 VDDHD VDDHD PCH L=60N W=1U M=2
MM8 CEBX BIST2 NET0284 VDDHD PCH L=60N W=500N M=1
MM10 NET0284 CEB VDDHD VDDHD PCH L=60N W=500N M=1
MM14 CEBX BIST1B NET0135 VDDHD PCH L=60N W=500N M=1
MN300 ENC EN VSSI VSSI NCH L=60N W=2U M=4
MM18 N7 CK1B NET0151 VSSI NCH L=60N W=1U M=1
MM11 NET0209 CEBM VSSI VSSI NCH L=60N W=500N M=1
MM17 CEBXL CEBX N7 VSSI NCH L=60N W=1U M=1
MM20 NET0151 RSC VSSI VSSI NCH L=60N W=1U M=2
MM3 CEBXL CK2 NET0168 VSSI NCH L=60N W=500N M=1
MM4 NET0168 EN NET0188 VSSI NCH L=60N W=500N M=1
MN200 ENC_Z EN VSSI VSSI NCH L=60N W=2U M=4
MM9 CEBX BIST1B NET0292 VSSI NCH L=60N W=500N M=1
MM5 NET0188 RSC VSSI VSSI NCH L=60N W=1U M=1
MN100 ENC_XY EN VSSI VSSI NCH L=60N W=2U M=4
MM13 CEBX BIST2 NET0209 VSSI NCH L=60N W=500N M=1
MM12 NET0292 CEB VSSI VSSI NCH L=60N W=500N M=1
XI141 CEBXL VSSI VDDHD EN S1AHSF400W40_AINV FN=2 WN=2U LN=0.06U FP=6 WP=1.4U LP=0.06U M=1
XI161 NET122 VSSI VDDHD EN_DCLK S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U 
+ LP=0.06U M=1
XI162 NET100 VSSI VDDHD NET0240 S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U 
+ LP=0.06U M=1
XINV5 NET0240 VSSI VDDHD NET94 S1AHSF400W40_AINV FN=3 WN=0.5U LN=0.06U FP=3 WP=1U 
+ LP=0.06U M=1
XI152 NET94 VSSI VDDHD EN_D S1AHSF400W40_AINV FN=6 WN=0.75U LN=0.06U FP=6 WP=1.6U 
+ LP=0.06U M=1
XINV10 NET112 VSSI VDDHD NET103 S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.3U 
+ LP=0.06U M=1
XINV8 NET115 VSSI VDDHD NET109 S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.3U 
+ LP=0.06U M=1
XINV9 NET109 VSSI VDDHD NET112 S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.3U 
+ LP=0.06U M=1
XINV7 EN VSSI VDDHD NET115 S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.3U LP=0.06U 
+ M=1
XI158 NET103 EN VSSI VDDHD NET100 S1AHSF400W40_ANOR FN2=1 WN2=0.3U LN2=0.06U FN1=1 
+ WN1=0.3U LN1=0.06U FP1=1 WP1=0.6U LP1=0.06U FP2=1 WP2=0.6U LP2=0.06U M=1
XNOR0 EN EN VSSI VDDHD NET122 S1AHSF400W40_ANOR FN2=1 WN2=0.3U LN2=0.06U FN1=1 WN1=0.3U 
+ LN1=0.06U FP1=1 WP1=0.6U LP1=0.06U FP2=1 WP2=0.6U LP2=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    ABUF_BIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ABUF_BIST A AM AX1B AX1BL AX1BL1B BIST1B BIST2 CK1B CK2 VDDHD VSSI
*.PININFO A:I AM:I BIST1B:I BIST2:I CK1B:I CK2:I AX1B:O AX1BL:O AX1BL1B:O 
*.PININFO VDDHD:B VSSI:B
MM24 AX BIST1B NET0124 VDDHD PCH L=60N W=600N M=1
MM25 NET0124 AM VDDHD VDDHD PCH L=60N W=600N M=1
MM26 AX1BL CK1B NET0149 VDDHD PCH L=60N W=300N M=1
MM27 NET0149 AX1BL1B VDDHD VDDHD PCH L=60N W=300N M=1
MM28 N5 CK2 VDDHD VDDHD PCH L=60N W=1U M=2
MM29 AX1BL AX1B N5 VDDHD PCH L=60N W=1U M=2
MM30 AX BIST2 NET0148 VDDHD PCH L=60N W=600N M=1
MM31 NET0148 A VDDHD VDDHD PCH L=60N W=600N M=1
MM16 AX BIST1B NET0113 VSSI NCH L=60N W=300N M=1
MM17 NET093 AM VSSI VSSI NCH L=60N W=300N M=1
MM18 AX BIST2 NET093 VSSI NCH L=60N W=300N M=1
MM19 AX1BL AX1B N7 VSSI NCH L=60N W=500N M=2
MM20 AX1BL CK2 NET078 VSSI NCH L=60N W=300N M=1
MM21 NET078 AX1BL1B VSSI VSSI NCH L=60N W=300N M=1
MM22 NET0113 A VSSI VSSI NCH L=60N W=300N M=1
MM23 N7 CK1B VSSI VSSI NCH L=60N W=500N M=2
XI39 AX VSSI VDDHD AX1B S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U LP=0.06U M=1
XI25 AX1BL VSSI VDDHD AX1BL1B S1AHSF400W40_AINV FN=2 WN=0.5U LN=0.06U FP=2 WP=1U LP=0.06U 
+ M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CDEC_BIST_M8M16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CDEC_BIST_M8M16 AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8] 
+ AX[9] AX[10] BIST1B BIST2 CEB CEBM CK1B CK2 CKP CKPD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] 
+ DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN ENC EN_DCLK PD REDEN REDENB 
+ RSC RW_RE VDDHD VDDI VSSI WEBXL WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] 
+ X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] 
+ XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO BIST1B:I BIST2:I CEB:I CEBM:I CKP:I CKPD:I CLK:I PD:I REDEN:I 
*.PININFO REDENB:I RSC:I WEBXL:I WEBXL1B:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I 
*.PININFO X[5]:I X[6]:I X[7]:I X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I 
*.PININFO XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I 
*.PININFO Y[0]:I Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AX[0]:O 
*.PININFO AX[1]:O AX[2]:O AX[3]:O AX[4]:O AX[5]:O AX[6]:O AX[7]:O AX[8]:O 
*.PININFO AX[9]:O AX[10]:O CK1B:O CK2:O DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O 
*.PININFO DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O 
*.PININFO DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O 
*.PININFO DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O 
*.PININFO DEC_X2[2]:O DEC_X2[3]:O DEC_X3[0]:O DEC_X3[1]:O DEC_X3[2]:O 
*.PININFO DEC_X3[3]:O DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O DEC_X3[7]:O 
*.PININFO DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O DEC_Y[5]:O 
*.PININFO DEC_Y[6]:O DEC_Y[7]:O EN:O ENC:O EN_DCLK:O RW_RE:O YL[0]:O VDDHD:B 
*.PININFO VDDI:B VSSI:B
XCEBBUF BIST1B BIST2 CEB CEBM CK1B CK2 EN ENC ENC_XY ENC_Z EN_D EN_DCLK RSC 
+ VDDHD VSSI S1AHSF400W40_ENBUFB_BIST
XABUF_Y<2> Y[2] YM[2] NET140 AYC[2] AYT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_X<3> X[3] XM[3] AX[3] AXC[3] AXT[3] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_X<4> X[4] XM[4] AX[4] AXC[4] AXT[4] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_X<5> X[5] XM[5] AX[5] AXC[5] AXT[5] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_X<8> X[8] XM[8] AX[8] AXC[8] AXT[8] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_X<9> X[9] XM[9] AX[9] AXC[9] AXT[9] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_X<10> X[10] XM[10] AX[10] AXC[10] AXT[10] BIST1B BIST2 CK1B CK2 VDDHD 
+ VSSI S1AHSF400W40_ABUF_BIST
XABUF_X<0> X[0] XM[0] AX[0] AXC[0] AXT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_X<1> X[1] XM[1] AX[1] AXC[1] AXT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_X<2> X[2] XM[2] AX[2] AXC[2] AXT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_Y<0> Y[0] YM[0] NET123[0] AYC[0] AYT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_Y<1> Y[1] YM[1] NET123[1] AYC[1] AYT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_X<6> X[6] XM[6] AX[6] AXC[6] AXT[6] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_X<7> X[7] XM[7] AX[7] AXC[7] AXT[7] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_Y<3> Y[3] YM[3] NET206 NET204 AYT[3] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XIDEC_YL CKPD CLK YL[0] EN_D ENC_XY AYT[3] VDDHD VSSI S1AHSF400W40_DECB1YL
XIPDEC_X0<0> AXC[0] AXT[0] AXC[1] AXT[1] AXC[2] XA[0] XA[1] XA[2] XA[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_X0<1> AXC[0] AXT[0] AXC[1] AXT[1] AXT[2] XA[4] XA[5] XA[6] XA[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_X3<0> AXC[8] AXT[8] AXC[9] AXT[9] AXC[10] Z[0] Z[1] Z[2] Z[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_X3<1> AXC[8] AXT[8] AXC[9] AXT[9] AXT[10] Z[4] Z[5] Z[6] Z[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_X1<0> AXC[3] AXT[3] AXC[4] AXT[4] AXC[5] XB[0] XB[1] XB[2] XB[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_X1<1> AXC[3] AXT[3] AXC[4] AXT[4] AXT[5] XB[4] XB[5] XB[6] XB[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_Y<0> AYC[0] AYT[0] AYC[1] AYT[1] AYC[2] XY[0] XY[1] XY[2] XY[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_Y<1> AYC[0] AYT[0] AYC[1] AYT[1] AYT[2] XY[4] XY[5] XY[6] XY[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIDEC_X0<0> CKPD CLK DEC_X0[0] EN_D ENC XA[0] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<1> CKPD CLK DEC_X0[1] EN_D ENC XA[1] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<2> CKPD CLK DEC_X0[2] EN_D ENC XA[2] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<3> CKPD CLK DEC_X0[3] EN_D ENC XA[3] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<4> CKPD CLK DEC_X0[4] EN_D ENC XA[4] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<5> CKPD CLK DEC_X0[5] EN_D ENC XA[5] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<6> CKPD CLK DEC_X0[6] EN_D ENC XA[6] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<7> CKPD CLK DEC_X0[7] EN_D ENC XA[7] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_RWRE CKPD CLK RW_RE EN_D ENC_XY WEBXL VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<0> CKPD CLK DEC_Y[0] EN_D ENC_XY XY[0] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<1> CKPD CLK DEC_Y[1] EN_D ENC_XY XY[1] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<2> CKPD CLK DEC_Y[2] EN_D ENC_XY XY[2] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<3> CKPD CLK DEC_Y[3] EN_D ENC_XY XY[3] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<0> CKP CLK DEC_X3[0] EN ENC_Z Z[0] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<1> CKP CLK DEC_X3[1] EN ENC_Z Z[1] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<2> CKP CLK DEC_X3[2] EN ENC_Z Z[2] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<3> CKP CLK DEC_X3[3] EN ENC_Z Z[3] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<4> CKP CLK DEC_X3[4] EN ENC_Z Z[4] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<5> CKP CLK DEC_X3[5] EN ENC_Z Z[5] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<6> CKP CLK DEC_X3[6] EN ENC_Z Z[6] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<7> CKP CLK DEC_X3[7] EN ENC_Z Z[7] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<4> CKPD CLK DEC_Y[4] EN_D ENC_XY XY[4] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<5> CKPD CLK DEC_Y[5] EN_D ENC_XY XY[5] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<6> CKPD CLK DEC_Y[6] EN_D ENC_XY XY[6] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<7> CKPD CLK DEC_Y[7] EN_D ENC_XY XY[7] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X2<0> CKPD CLK DEC_X2[0] EN_D ENC_XY XC[0] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X2<1> CKPD CLK DEC_X2[1] EN_D ENC_XY XC[1] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X2<2> CKPD CLK DEC_X2[2] EN_D ENC_XY XC[2] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X2<3> CKPD CLK DEC_X2[3] EN_D ENC_XY XC[3] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<0> CKPD CLK DEC_X1[0] EN_D ENC XB[0] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<1> CKPD CLK DEC_X1[1] EN_D ENC XB[1] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<2> CKPD CLK DEC_X1[2] EN_D ENC XB[2] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<3> CKPD CLK DEC_X1[3] EN_D ENC XB[3] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<4> CKPD CLK DEC_X1[4] EN_D ENC XB[4] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<5> CKPD CLK DEC_X1[5] EN_D ENC XB[5] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<6> CKPD CLK DEC_X1[6] EN_D ENC XB[6] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<7> CKPD CLK DEC_X1[7] EN_D ENC XB[7] VDDHD VSSI S1AHSF400W40_DECB1
XIPDEC_X2<0> AXC[6] AXT[6] AXC[7] XC[0] XC[1] VDDHD VSSI S1AHSF400W40_DECB2
XIPDEC_X2<1> AXC[6] AXT[6] AXT[7] XC[2] XC[3] VDDHD VSSI S1AHSF400W40_DECB2
XCKBUF CK1B CK2 CKPD CLK VDDHD VSSI S1AHSF400W40_CKBUF
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_F_M16_BIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_F_M16_BIST AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD 
+ PD_BUF PD_CVDDBUF PTSEL REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL 
+ VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] 
+ WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] 
+ XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] 
+ Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I REDEN:I REDENB:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I 
*.PININFO XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I 
*.PININFO Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O BIST2IO:O 
*.PININFO BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O 
*.PININFO DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O DEC_X1[0]:O 
*.PININFO DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O DEC_X1[5]:O 
*.PININFO DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O DEC_X2[2]:O 
*.PININFO DEC_X2[3]:O DEC_X3[0]:O DEC_X3[1]:O DEC_X3[2]:O DEC_X3[3]:O 
*.PININFO DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O DEC_X3[7]:O DEC_Y[0]:O 
*.PININFO DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O 
*.PININFO DEC_Y[7]:O PD_BUF:O PD_CVDDBUF:O RW_RE:O VHI:O VLO:O WLP_SAE:O 
*.PININFO WLP_SAEB:O YL[0]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE_TK:B
XCOTHERS AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKD CKP CKPD 
+ CLK EN ENC EN_DCLK PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WEB WEBM WEBXL WEBXL1B WLP_SAE WLP_SAEB WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2] S1AHSF400W40_COTH_F_BIST
XCDEC AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8] AX[9] AX[10] 
+ BIST1B BIST2 CEB CEBM CK1B CK2 CKP CKPD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN ENC EN_DCLK PD REDEN REDENB RSC RW_RE 
+ VDDHD VDDI VSSI WEBXL WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] 
+ X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] 
+ XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3] S1AHSF400W40_CDEC_BIST_M8M16
MX0_PD<0> DEC_X0[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<1> DEC_X0[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<2> DEC_X0[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<3> DEC_X0[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<4> DEC_X0[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<5> DEC_X0[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<6> DEC_X0[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<7> DEC_X0[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<0> DEC_X1[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<1> DEC_X1[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<2> DEC_X1[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<3> DEC_X1[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<4> DEC_X1[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<5> DEC_X1[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<6> DEC_X1[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<7> DEC_X1[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_F_M8_BIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_F_M8_BIST AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD 
+ PD_BUF PD_CVDDBUF PTSEL REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL 
+ VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] 
+ WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] 
+ XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] 
+ Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I REDEN:I REDENB:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I 
*.PININFO XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I 
*.PININFO Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O BIST2IO:O 
*.PININFO BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O 
*.PININFO DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O DEC_X1[0]:O 
*.PININFO DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O DEC_X1[5]:O 
*.PININFO DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O DEC_X2[2]:O 
*.PININFO DEC_X2[3]:O DEC_X3[0]:O DEC_X3[1]:O DEC_X3[2]:O DEC_X3[3]:O 
*.PININFO DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O DEC_X3[7]:O DEC_Y[0]:O 
*.PININFO DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O 
*.PININFO DEC_Y[7]:O PD_BUF:O PD_CVDDBUF:O RW_RE:O VHI:O VLO:O WLP_SAE:O 
*.PININFO WLP_SAEB:O YL[0]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE_TK:B
XCOTHERS AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKD CKP CKPD 
+ CLK EN ENC EN_DCLK PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WEB WEBM WEBXL WEBXL1B WLP_SAE WLP_SAEB WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2] S1AHSF400W40_COTH_F_BIST
XCDEC AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8] AX[9] AX[10] 
+ BIST1B BIST2 CEB CEBM CK1B CK2 CKP CKPD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN ENC EN_DCLK PD REDEN REDENB RSC RW_RE 
+ VDDHD VDDI VSSI WEBXL WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] 
+ X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] 
+ XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3] S1AHSF400W40_CDEC_BIST_M8M16
MX0_PD<0> DEC_X0[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<1> DEC_X0[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<2> DEC_X0[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<3> DEC_X0[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<4> DEC_X0[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<5> DEC_X0[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<6> DEC_X0[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<7> DEC_X0[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<0> DEC_X1[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<1> DEC_X1[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<2> DEC_X1[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<3> DEC_X1[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<4> DEC_X1[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<5> DEC_X1[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<6> DEC_X1[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<7> DEC_X1[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CDEC_BIST_M4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CDEC_BIST_M4 AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8] 
+ AX[9] AX[10] BIST1B BIST2 CEB CEBM CK1B CK2 CKP CKPD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] 
+ DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN ENC EN_DCLK PD REDEN REDENB 
+ RSC RW_RE VDDHD VDDI VSSI WEBXL WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] 
+ X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] 
+ XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO BIST1B:I BIST2:I CEB:I CEBM:I CKP:I CKPD:I CLK:I PD:I REDEN:I 
*.PININFO REDENB:I RSC:I WEBXL:I WEBXL1B:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I 
*.PININFO X[5]:I X[6]:I X[7]:I X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I 
*.PININFO XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I 
*.PININFO Y[0]:I Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AX[0]:O 
*.PININFO AX[1]:O AX[2]:O AX[3]:O AX[4]:O AX[5]:O AX[6]:O AX[7]:O AX[8]:O 
*.PININFO AX[9]:O AX[10]:O CK1B:O CK2:O DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O 
*.PININFO DEC_X0[3]:O DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O 
*.PININFO DEC_X1[0]:O DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O 
*.PININFO DEC_X1[5]:O DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O 
*.PININFO DEC_X2[2]:O DEC_X2[3]:O DEC_X3[0]:O DEC_X3[1]:O DEC_X3[2]:O 
*.PININFO DEC_X3[3]:O DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O DEC_X3[7]:O 
*.PININFO DEC_Y[0]:O DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O DEC_Y[5]:O 
*.PININFO DEC_Y[6]:O DEC_Y[7]:O EN:O ENC:O EN_DCLK:O RW_RE:O YL[0]:O VDDHD:B 
*.PININFO VDDI:B VSSI:B
XCEBBUF BIST1B BIST2 CEB CEBM CK1B CK2 EN ENC ENC_XY ENC_Z EN_D EN_DCLK RSC 
+ VDDHD VSSI S1AHSF400W40_ENBUFB_BIST
XABUF_X<6> X[6] XM[6] AX[6] AXC[6] AXT[6] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_X<7> X[7] XM[7] AX[7] AXC[7] AXT[7] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_Y<3> Y[3] YM[3] NET0283 NET207 AYT[3] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_Y<2> Y[2] YM[2] NET0294 NET217 NET216 BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_X<3> X[3] XM[3] AX[3] AXC[3] AXT[3] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_X<4> X[4] XM[4] AX[4] AXC[4] AXT[4] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_X<5> X[5] XM[5] AX[5] AXC[5] AXT[5] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_X<8> X[8] XM[8] AX[8] AXC[8] AXT[8] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_X<9> X[9] XM[9] AX[9] AXC[9] AXT[9] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_X<10> X[10] XM[10] AX[10] AXC[10] AXT[10] BIST1B BIST2 CK1B CK2 VDDHD 
+ VSSI S1AHSF400W40_ABUF_BIST
XABUF_X<0> X[0] XM[0] AX[0] AXC[0] AXT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_X<1> X[1] XM[1] AX[1] AXC[1] AXT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_X<2> X[2] XM[2] AX[2] AXC[2] AXT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_Y<0> Y[0] YM[0] NET089[0] AYC[0] AYT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XABUF_Y<1> Y[1] YM[1] NET089[1] AYC[1] AYT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST
XIDEC_YL CKPD CLK YL[0] EN_D ENC_XY AYT[3] VDDHD VSSI S1AHSF400W40_DECB1YL
XCKBUF CK1B CK2 CKPD CLK VDDHD VSSI S1AHSF400W40_CKBUF
XIPDEC_X2<0> AXC[6] AXT[6] AXC[7] XC[0] XC[1] VDDHD VSSI S1AHSF400W40_DECB2
XIPDEC_X2<1> AXC[6] AXT[6] AXT[7] XC[2] XC[3] VDDHD VSSI S1AHSF400W40_DECB2
XIDEC_X3<0> CKP CLK DEC_X3[0] EN ENC_Z Z[0] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<1> CKP CLK DEC_X3[1] EN ENC_Z Z[1] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<2> CKP CLK DEC_X3[2] EN ENC_Z Z[2] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<3> CKP CLK DEC_X3[3] EN ENC_Z Z[3] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<4> CKP CLK DEC_X3[4] EN ENC_Z Z[4] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<5> CKP CLK DEC_X3[5] EN ENC_Z Z[5] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<6> CKP CLK DEC_X3[6] EN ENC_Z Z[6] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X3<7> CKP CLK DEC_X3[7] EN ENC_Z Z[7] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X2<0> CKPD CLK DEC_X2[0] EN_D ENC_XY XC[0] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X2<1> CKPD CLK DEC_X2[1] EN_D ENC_XY XC[1] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X2<2> CKPD CLK DEC_X2[2] EN_D ENC_XY XC[2] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X2<3> CKPD CLK DEC_X2[3] EN_D ENC_XY XC[3] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<0> CKPD CLK DEC_X1[0] EN_D ENC XB[0] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<1> CKPD CLK DEC_X1[1] EN_D ENC XB[1] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<2> CKPD CLK DEC_X1[2] EN_D ENC XB[2] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<3> CKPD CLK DEC_X1[3] EN_D ENC XB[3] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<4> CKPD CLK DEC_X1[4] EN_D ENC XB[4] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<5> CKPD CLK DEC_X1[5] EN_D ENC XB[5] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<6> CKPD CLK DEC_X1[6] EN_D ENC XB[6] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X1<7> CKPD CLK DEC_X1[7] EN_D ENC XB[7] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<0> CKPD CLK DEC_X0[0] EN_D ENC XA[0] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<1> CKPD CLK DEC_X0[1] EN_D ENC XA[1] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<2> CKPD CLK DEC_X0[2] EN_D ENC XA[2] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<3> CKPD CLK DEC_X0[3] EN_D ENC XA[3] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<4> CKPD CLK DEC_X0[4] EN_D ENC XA[4] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<5> CKPD CLK DEC_X0[5] EN_D ENC XA[5] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<6> CKPD CLK DEC_X0[6] EN_D ENC XA[6] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_X0<7> CKPD CLK DEC_X0[7] EN_D ENC XA[7] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_RWRE CKPD CLK RW_RE EN_D ENC_XY WEBXL VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<4> CKPD CLK DEC_Y[4] EN_D ENC_XY XY[4] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<5> CKPD CLK DEC_Y[5] EN_D ENC_XY XY[5] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<6> CKPD CLK DEC_Y[6] EN_D ENC_XY XY[6] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<7> CKPD CLK DEC_Y[7] EN_D ENC_XY XY[7] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<0> CKPD CLK DEC_Y[0] EN_D ENC_XY XY[0] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<1> CKPD CLK DEC_Y[1] EN_D ENC_XY XY[1] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<2> CKPD CLK DEC_Y[2] EN_D ENC_XY XY[2] VDDHD VSSI S1AHSF400W40_DECB1
XIDEC_Y<3> CKPD CLK DEC_Y[3] EN_D ENC_XY XY[3] VDDHD VSSI S1AHSF400W40_DECB1
XIPDEC_X0<0> AXC[0] AXT[0] AXC[1] AXT[1] AXC[2] XA[0] XA[1] XA[2] XA[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_X0<1> AXC[0] AXT[0] AXC[1] AXT[1] AXT[2] XA[4] XA[5] XA[6] XA[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_Y<0> AYC[0] AYT[0] AYC[1] AYT[1] WEBXL XY[0] XY[1] XY[2] XY[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_Y<1> AYC[0] AYT[0] AYC[1] AYT[1] WEBXL1B XY[4] XY[5] XY[6] XY[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_X3<0> AXC[8] AXT[8] AXC[9] AXT[9] AXC[10] Z[0] Z[1] Z[2] Z[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_X3<1> AXC[8] AXT[8] AXC[9] AXT[9] AXT[10] Z[4] Z[5] Z[6] Z[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_X1<0> AXC[3] AXT[3] AXC[4] AXT[4] AXC[5] XB[0] XB[1] XB[2] XB[3] VDDHD 
+ VSSI S1AHSF400W40_DECB4
XIPDEC_X1<1> AXC[3] AXT[3] AXC[4] AXT[4] AXT[5] XB[4] XB[5] XB[6] XB[7] VDDHD 
+ VSSI S1AHSF400W40_DECB4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_F_M4_BIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_F_M4_BIST AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD 
+ PD_BUF PD_CVDDBUF PTSEL REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL 
+ VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] 
+ WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] 
+ XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] 
+ Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I REDEN:I REDENB:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I 
*.PININFO XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I 
*.PININFO Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O BIST2IO:O 
*.PININFO BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O 
*.PININFO DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O DEC_X1[0]:O 
*.PININFO DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O DEC_X1[5]:O 
*.PININFO DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O DEC_X2[2]:O 
*.PININFO DEC_X2[3]:O DEC_X3[0]:O DEC_X3[1]:O DEC_X3[2]:O DEC_X3[3]:O 
*.PININFO DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O DEC_X3[7]:O DEC_Y[0]:O 
*.PININFO DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O 
*.PININFO DEC_Y[7]:O PD_BUF:O PD_CVDDBUF:O RW_RE:O VHI:O VLO:O WLP_SAE:O 
*.PININFO WLP_SAEB:O YL[0]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE_TK:B
XCOTHERS AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKD CKP CKPD 
+ CLK EN ENC EN_DCLK PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WEB WEBM WEBXL WEBXL1B WLP_SAE WLP_SAEB WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2] S1AHSF400W40_COTH_F_BIST
XCDEC AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8] AX[9] AX[10] 
+ BIST1B BIST2 CEB CEBM CK1B CK2 CKP CKPD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN ENC EN_DCLK PD REDEN REDENB RSC RW_RE 
+ VDDHD VDDI VSSI WEBXL WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] 
+ X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] 
+ XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3] S1AHSF400W40_CDEC_BIST_M4
MX0_PD<0> DEC_X0[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<1> DEC_X0[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<2> DEC_X0[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<3> DEC_X0[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<4> DEC_X0[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<5> DEC_X0[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<6> DEC_X0[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<7> DEC_X0[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<0> DEC_X1[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<1> DEC_X1[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<2> DEC_X1[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<3> DEC_X1[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<4> DEC_X1[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<5> DEC_X1[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<6> DEC_X1[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<7> DEC_X1[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    RESETD
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_RESETD BLTRKWLDRV CK2 CKP CKPD CKPDCLK IOSAEB RSTCK TK TRKBL VDDHD 
+ VSSI WEBXL WLP_SAE WLP_SAE_TK PTSEL RV[0] RV[1] WV[0] WV[1] WV[2]
*.PININFO CK2:I CKP:I WEBXL:I PTSEL:I RV[0]:I RV[1]:I WV[0]:I WV[1]:I WV[2]:I 
*.PININFO BLTRKWLDRV:O CKPD:O CKPDCLK:O IOSAEB:O RSTCK:O WLP_SAE:O TK:B 
*.PININFO TRKBL:B VDDHD:B VSSI:B WLP_SAE_TK:B
XTSEL_READ CKP RV[0] RV[1] VDDHD VSSI RTD_01_11 RTD_10 S1AHSF400W40_RESETD_TSEL
XI616 TRKBL3B WV[0] WV[1] VDDHD VSSI WTD_01_11 WTD_10 S1AHSF400W40_RESETD_TSEL
MP16 WLP_SAE NET0346 VDDHD VDDHD PCH L=60N W=2U M=6
MN7 WLP_SAE NET0346 VSSI VSSI NCH L=60N W=1U M=6
XI584 CKP RTD_01_11 RTD_10 VSSI VDDHD RTKB S1AHSF400W40_ANAND3 FN3=1 WN3=1.2U LN3=60N 
+ FN2=1 WN2=1.2U LN2=60N FN1=1 WN1=1.2U LN1=60N FP1=1 WP1=0.8U LP1=60N FP2=1 
+ WP2=0.8U LP2=60N FP3=1 WP3=0.8U LP3=60N M=1
XI612 TRKBL3B WTD_01_11 WTD_10 VSSI VDDHD NET0346 S1AHSF400W40_ANAND3 FN3=2 WN3=1.5U 
+ LN3=60N FN2=2 WN2=1.5U LN2=60N FN1=2 WN1=1.5U LN1=60N FP1=2 WP1=1U LP1=60N 
+ FP2=2 WP2=1U LP2=60N FP3=2 WP3=1U LP3=60N M=1
XNAND4 TRKBL1B CKP VSSI VDDHD RSTCKB S1AHSF400W40_ANAND FN2=1 WN2=0.8U LN2=0.06U FN1=1 
+ WN1=0.8U LN1=0.06U FP1=1 WP1=0.6U LP1=0.06U FP2=1 WP2=0.6U LP2=0.06U M=1
XI592 Z6 Z5 VSSI VDDHD Z7 S1AHSF400W40_ANAND FN2=1 WN2=0.25U LN2=0.06U FN1=1 WN1=0.25U 
+ LN1=0.06U FP1=1 WP1=0.3U LP1=0.06U FP2=1 WP2=0.3U LP2=0.06U M=1
XI521 WLP_SAE3B WLP_SAE_TK1B VSSI VDDHD NET342 S1AHSF400W40_ANAND FN2=1 WN2=0.25U 
+ LN2=0.06U FN1=1 WN1=0.25U LN1=0.06U FP1=1 WP1=0.3U LP1=0.06U FP2=1 WP2=0.3U 
+ LP2=0.06U M=1
XI575 WEBXL TRKBL1B VSSI VDDHD TRKBL2 S1AHSF400W40_ANAND FN2=1 WN2=0.8U LN2=60N FN1=1 
+ WN1=0.8U LN1=60N FP1=1 WP1=0.6U LP1=60N FP2=1 WP2=0.6U LP2=60N M=1
XI589 Z3 VSSI VDDHD Z4 S1AHSF400W40_AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=0.4U LP=0.06U M=1
XI598 WLP_SAE VSSI VDDHD WLP_SAE_1B S1AHSF400W40_AINV FN=1 WN=0.4U LN=0.06U FP=1 WP=0.4U 
+ LP=0.06U M=1
XI601 WLP_SAE2 VSSI VDDHD WLP_SAE3B S1AHSF400W40_AINV FN=1 WN=0.4U LN=0.06U FP=1 WP=0.4U 
+ LP=0.06U M=1
XI620 RSTCKB VSSI VDDHD RSTCK S1AHSF400W40_AINV FN=1 WN=0.4U LN=60N FP=1 WP=0.6U LP=60N 
+ M=2
XI618 NET327 VSSI VDDHD NET299 S1AHSF400W40_AINV FN=2 WN=0.75U LN=60N FP=2 WP=1.5U LP=60N 
+ M=1
*XI585 Z0 VSSI VDDHD Z1 AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=0.4U LP=0.06U M=1
XI586 Z6 VSSI VDDHD Z0 S1AHSF400W40_AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=0.4U LP=0.06U M=1
XI606 CKPD VSSI VDDHD Z10 S1AHSF400W40_AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=0.4U LP=0.06U 
+ M=1
XI607 Z10 VSSI VDDHD CKPDCLK S1AHSF400W40_AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=0.4U 
+ LP=0.06U M=1
XI594 Z8 VSSI VDDHD CKPD S1AHSF400W40_AINV FN=8 WN=0.3U LN=0.06U FP=8 WP=0.6U LP=0.06U M=1
XI593 Z7 VSSI VDDHD Z8 S1AHSF400W40_AINV FN=2 WN=0.3U LN=0.06U FP=2 WP=0.6U LP=0.06U M=1
XI566 WLP_SAE_TK VSSI VDDHD WLP_SAE_TK1B S1AHSF400W40_AINV FN=1 WN=0.4U LN=0.06U FP=1 
+ WP=0.4U LP=0.06U M=1
XI600 WLP_SAE_1B VSSI VDDHD WLP_SAE2 S1AHSF400W40_AINV FN=1 WN=0.4U LN=0.06U FP=1 WP=0.4U 
+ LP=0.06U M=1
XI591 CKP VSSI VDDHD Z6 S1AHSF400W40_AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=0.4U LP=0.06U M=1
XI619 NET342 VSSI VDDHD NET327 S1AHSF400W40_AINV FN=1 WN=0.4U LN=60N FP=1 WP=0.8U LP=60N 
+ M=1
XI617 NET299 VSSI VDDHD IOSAEB S1AHSF400W40_AINV FN=8 WN=0.75U LN=60N FP=8 WP=1.5U LP=60N 
+ M=1
XI537 RTKB2 VSSI VDDHD BLTRKWLDRV S1AHSF400W40_AINV FN=8 WN=0.75U LN=60N FP=8 WP=1.5U 
+ LP=60N M=1
XI613 TRKBL2 VSSI VDDHD TRKBL3B S1AHSF400W40_AINV FN=1 WN=0.4U LN=0.06U FP=1 WP=0.6U 
+ LP=0.06U M=1
XI588 Z0 VSSI VDDHD Z3 S1AHSF400W40_AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=0.4U LP=0.06U M=1
XI590 Z4 VSSI VDDHD Z5 S1AHSF400W40_AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=0.4U LP=0.06U M=1
XI541 RTKB VSSI VDDHD RTKB1B S1AHSF400W40_AINV FN=1 WN=0.4U LN=60N FP=1 WP=0.8U LP=60N M=1
XI574 TRKBL VSSI VDDHD TRKBL1B S1AHSF400W40_AINV FN=1 WN=0.4U LN=60N FP=1 WP=0.8U LP=60N 
+ M=1
XI540 RTKB1B VSSI VDDHD RTKB2 S1AHSF400W40_AINV FN=2 WN=0.75U LN=60N FP=2 WP=1.5U LP=60N 
+ M=1
*XI587 Z1 VSSI VDDHD Z2 AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=0.4U LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    COTH_BIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_COTH_BIST AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKD 
+ CKP CKPD CLK EN ENC_D EN_D PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL 
+ VDDHD VDDI VHI VLO VSSI WEB WEBM WEBXL WEBXL1B WLP_SAE WLP_SAEB WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2]
*.PININFO AWT:I BIST:I CK1B:I CK2:I CLK:I EN:I ENC_D:I EN_D:I PD:I PTSEL:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I AWT2:O BIST1B:O BIST2:O BIST2IO:O BLTRKWLDRV:O CKD:O 
*.PININFO CKP:O CKPD:O PD_BUF:O RSC:O VHI:O VLO:O WEBXL:O WEBXL1B:O WLP_SAE:O 
*.PININFO WLP_SAEB:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE_TK:B
XVHILO_SB VDDHD VHI VLO VSSI S1AHSF400W40_VHILO_SB
XWEBBUF BIST1B BIST2 CK1B CK2 VDDHD VSSI WEB WEBM WEBXL WEBXL1B S1AHSF400W40_WEBBUF_BIST
XIDEC_CKD CKPDCLK CLK CKD EN_D ENC_D WEBXL1B VDDHD VSSI S1AHSF400W40_DECB1
XAWTD AWT AWT2 PD VDDHD VDDI VSSI S1AHSF400W40_AWTD
XBISTD BIST BIST1B BIST2 BIST2IO VDDHD VSSI S1AHSF400W40_BISTD
XCKG CKP CLK EN RSC RSTCK TM VDDHD VSSI S1AHSF400W40_CKG
XRESETD BLTRKWLDRV CK2 CKP CKPD CKPDCLK WLP_SAEB RSTCK TK TRKBL VDDHD VSSI 
+ WEBXL WLP_SAE WLP_SAE_TK PTSEL RTSEL[0] RTSEL[1] WTSEL[0] WTSEL[1] WTSEL[2] 
+ S1AHSF400W40_RESETD
XPDBUF PD PD_BUF VDDI VSSI S1AHSF400W40_PDBUF
MP2 VDDHD PD VDDI VDDI PCH L=60N W=5U M=19
MP1 VDDHD PD VDDI VDDI PCH L=60N W=3.5U M=8
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_M16_BIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_M16_BIST AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD 
+ PD_BUF PD_CVDDBUF PTSEL REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL 
+ VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] 
+ WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] 
+ XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] 
+ Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I REDEN:I REDENB:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I 
*.PININFO XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I 
*.PININFO Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O BIST2IO:O 
*.PININFO BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O 
*.PININFO DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O DEC_X1[0]:O 
*.PININFO DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O DEC_X1[5]:O 
*.PININFO DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O DEC_X2[2]:O 
*.PININFO DEC_X2[3]:O DEC_X3[0]:O DEC_X3[1]:O DEC_X3[2]:O DEC_X3[3]:O 
*.PININFO DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O DEC_X3[7]:O DEC_Y[0]:O 
*.PININFO DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O 
*.PININFO DEC_Y[7]:O PD_BUF:O PD_CVDDBUF:O RW_RE:O VHI:O VLO:O WLP_SAE:O 
*.PININFO WLP_SAEB:O YL[0]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE_TK:B
XCOTHERS AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKD CKP CKPD 
+ CLK EN ENC EN_DCLK PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WEB WEBM WEBXL WEBXL1B WLP_SAE WLP_SAEB WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2] S1AHSF400W40_COTH_BIST
XCDEC AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8] AX[9] AX[10] 
+ BIST1B BIST2 CEB CEBM CK1B CK2 CKP CKPD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN ENC EN_DCLK PD REDEN REDENB RSC RW_RE 
+ VDDHD VDDI VSSI WEBXL WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] 
+ X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] 
+ XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3] S1AHSF400W40_CDEC_BIST_M8M16
MX0_PD<0> DEC_X0[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<1> DEC_X0[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<2> DEC_X0[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<3> DEC_X0[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<4> DEC_X0[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<5> DEC_X0[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<6> DEC_X0[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<7> DEC_X0[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<0> DEC_X1[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<1> DEC_X1[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<2> DEC_X1[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<3> DEC_X1[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<4> DEC_X1[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<5> DEC_X1[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<6> DEC_X1[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<7> DEC_X1[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_M8_BIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_M8_BIST AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD 
+ PD_BUF PD_CVDDBUF PTSEL REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL 
+ VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] 
+ WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] 
+ XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] 
+ Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I REDEN:I REDENB:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I 
*.PININFO XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I 
*.PININFO Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O BIST2IO:O 
*.PININFO BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O 
*.PININFO DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O DEC_X1[0]:O 
*.PININFO DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O DEC_X1[5]:O 
*.PININFO DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O DEC_X2[2]:O 
*.PININFO DEC_X2[3]:O DEC_X3[0]:O DEC_X3[1]:O DEC_X3[2]:O DEC_X3[3]:O 
*.PININFO DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O DEC_X3[7]:O DEC_Y[0]:O 
*.PININFO DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O 
*.PININFO DEC_Y[7]:O PD_BUF:O PD_CVDDBUF:O RW_RE:O VHI:O VLO:O WLP_SAE:O 
*.PININFO WLP_SAEB:O YL[0]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE_TK:B
XCOTHERS AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKD CKP CKPD 
+ CLK EN ENC EN_DCLK PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WEB WEBM WEBXL WEBXL1B WLP_SAE WLP_SAEB WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2] S1AHSF400W40_COTH_BIST
XCDEC AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8] AX[9] AX[10] 
+ BIST1B BIST2 CEB CEBM CK1B CK2 CKP CKPD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN ENC EN_DCLK PD REDEN REDENB RSC RW_RE 
+ VDDHD VDDI VSSI WEBXL WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] 
+ X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] 
+ XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3] S1AHSF400W40_CDEC_BIST_M8M16
MX0_PD<0> DEC_X0[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<1> DEC_X0[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<2> DEC_X0[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<3> DEC_X0[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<4> DEC_X0[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<5> DEC_X0[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<6> DEC_X0[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<7> DEC_X0[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<0> DEC_X1[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<1> DEC_X1[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<2> DEC_X1[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<3> DEC_X1[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<4> DEC_X1[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<5> DEC_X1[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<6> DEC_X1[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<7> DEC_X1[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_M4_BIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_M4_BIST AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD 
+ PD_BUF PD_CVDDBUF PTSEL REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL 
+ VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] 
+ WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] 
+ XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] 
+ Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I REDEN:I REDENB:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I 
*.PININFO XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I 
*.PININFO Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O BIST2IO:O 
*.PININFO BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O 
*.PININFO DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O DEC_X1[0]:O 
*.PININFO DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O DEC_X1[5]:O 
*.PININFO DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O DEC_X2[2]:O 
*.PININFO DEC_X2[3]:O DEC_X3[0]:O DEC_X3[1]:O DEC_X3[2]:O DEC_X3[3]:O 
*.PININFO DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O DEC_X3[7]:O DEC_Y[0]:O 
*.PININFO DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O 
*.PININFO DEC_Y[7]:O PD_BUF:O PD_CVDDBUF:O RW_RE:O VHI:O VLO:O WLP_SAE:O 
*.PININFO WLP_SAEB:O YL[0]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE_TK:B
XCOTHERS AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKD CKP CKPD 
+ CLK EN ENC EN_DCLK PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WEB WEBM WEBXL WEBXL1B WLP_SAE WLP_SAEB WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2] S1AHSF400W40_COTH_BIST
XCDEC AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8] AX[9] AX[10] 
+ BIST1B BIST2 CEB CEBM CK1B CK2 CKP CKPD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN ENC EN_DCLK PD REDEN REDENB RSC RW_RE 
+ VDDHD VDDI VSSI WEBXL WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] 
+ X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] 
+ XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3] S1AHSF400W40_CDEC_BIST_M4
MX0_PD<0> DEC_X0[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<1> DEC_X0[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<2> DEC_X0[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<3> DEC_X0[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<4> DEC_X0[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<5> DEC_X0[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<6> DEC_X0[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<7> DEC_X0[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<0> DEC_X1[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<1> DEC_X1[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<2> DEC_X1[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<3> DEC_X1[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<4> DEC_X1[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<5> DEC_X1[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<6> DEC_X1[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<7> DEC_X1[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    COTH
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_COTH AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKD CKP 
+ CKPD CLK EN ENC_D EN_D PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL 
+ VDDHD VDDI VHI VLO VSSI WEB WEBM WEBXL WEBXL1B WLP_SAE WLP_SAEB WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2]
*.PININFO AWT:I BIST:I CK1B:I CK2:I CLK:I EN:I ENC_D:I EN_D:I PD:I PTSEL:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I AWT2:O BIST1B:O BIST2:O BIST2IO:O BLTRKWLDRV:O CKD:O 
*.PININFO CKP:O CKPD:O PD_BUF:O RSC:O VHI:O VLO:O WEBXL:O WEBXL1B:O WLP_SAE:O 
*.PININFO WLP_SAEB:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE_TK:B
XRESETD BLTRKWLDRV CK2 CKP CKPD CKPDCLK WLP_SAEB RSTCK TK TRKBL VDDHD VSSI 
+ WEBXL WLP_SAE WLP_SAE_TK PTSEL RTSEL[0] RTSEL[1] WTSEL[0] WTSEL[1] WTSEL[2] 
+ S1AHSF400W40_RESETD
XIDEC_CKD CKPDCLK CLK CKD EN_D ENC_D WEBXL1B VDDHD VSSI S1AHSF400W40_DECB1
XWEBBUF BIST1B BIST2 CK1B CK2 VDDHD VSSI WEB WEBM WEBXL WEBXL1B S1AHSF400W40_WEBBUF
XVHILO VDDHD VHI VLO VSSI S1AHSF400W40_VHILO
XAWTD AWT AWT2 PD VDDHD VDDI VSSI S1AHSF400W40_AWTD
XBISTD BIST BIST1B BIST2 BIST2IO VDDHD VSSI S1AHSF400W40_BISTD
XCKG CKP CLK EN RSC RSTCK TM VDDHD VSSI S1AHSF400W40_CKG
XPDBUF PD PD_BUF VDDI VSSI S1AHSF400W40_PDBUF
MP2 VDDHD PD VDDI VDDI PCH L=60N W=5U M=19
MP1 VDDHD PD VDDI VDDI PCH L=60N W=3.5U M=8
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_M4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_M4 AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD 
+ PD_BUF PD_CVDDBUF PTSEL REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL 
+ VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] 
+ WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] 
+ XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] 
+ Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I REDEN:I REDENB:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I 
*.PININFO XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I 
*.PININFO Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O BIST2IO:O 
*.PININFO BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O 
*.PININFO DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O DEC_X1[0]:O 
*.PININFO DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O DEC_X1[5]:O 
*.PININFO DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O DEC_X2[2]:O 
*.PININFO DEC_X2[3]:O DEC_X3[0]:O DEC_X3[1]:O DEC_X3[2]:O DEC_X3[3]:O 
*.PININFO DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O DEC_X3[7]:O DEC_Y[0]:O 
*.PININFO DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O 
*.PININFO DEC_Y[7]:O PD_BUF:O PD_CVDDBUF:O RW_RE:O VHI:O VLO:O WLP_SAE:O 
*.PININFO WLP_SAEB:O YL[0]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE_TK:B
MX0_PD<0> DEC_X0[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<1> DEC_X0[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<2> DEC_X0[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<3> DEC_X0[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<4> DEC_X0[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<5> DEC_X0[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<6> DEC_X0[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<7> DEC_X0[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<0> DEC_X1[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<1> DEC_X1[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<2> DEC_X1[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<3> DEC_X1[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<4> DEC_X1[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<5> DEC_X1[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<6> DEC_X1[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<7> DEC_X1[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
XCOTHERS AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKD CKP CKPD 
+ CLK EN ENC EN_DCLK PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WEB WEBM WEBXL WEBXL1B WLP_SAE WLP_SAEB WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2] S1AHSF400W40_COTH
XCDEC AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8] AX[9] AX[10] 
+ BIST1B BIST2 CEB CEBM CK1B CK2 CKP CKPD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN ENC EN_DCLK PD REDEN REDENB RSC RW_RE 
+ VDDHD VDDI VSSI WEBXL WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] 
+ X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] 
+ XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3] S1AHSF400W40_CDEC_M4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_M16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_M16 AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD 
+ PD_BUF PD_CVDDBUF PTSEL REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL 
+ VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] 
+ WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] 
+ XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] 
+ Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I REDEN:I REDENB:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I 
*.PININFO XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I 
*.PININFO Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O BIST2IO:O 
*.PININFO BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O 
*.PININFO DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O DEC_X1[0]:O 
*.PININFO DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O DEC_X1[5]:O 
*.PININFO DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O DEC_X2[2]:O 
*.PININFO DEC_X2[3]:O DEC_X3[0]:O DEC_X3[1]:O DEC_X3[2]:O DEC_X3[3]:O 
*.PININFO DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O DEC_X3[7]:O DEC_Y[0]:O 
*.PININFO DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O 
*.PININFO DEC_Y[7]:O PD_BUF:O PD_CVDDBUF:O RW_RE:O VHI:O VLO:O WLP_SAE:O 
*.PININFO WLP_SAEB:O YL[0]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE_TK:B
XCOTHERS AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKD CKP CKPD 
+ CLK EN ENC EN_DCLK PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WEB WEBM WEBXL WEBXL1B WLP_SAE WLP_SAEB WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2] S1AHSF400W40_COTH
XCDEC AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8] AX[9] AX[10] 
+ BIST1B BIST2 CEB CEBM CK1B CK2 CKP CKPD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN ENC EN_DCLK PD REDEN REDENB RSC RW_RE 
+ VDDHD VDDI VSSI WEBXL WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] 
+ X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] 
+ XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3] S1AHSF400W40_CDEC_M8M16
MX0_PD<0> DEC_X0[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<1> DEC_X0[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<2> DEC_X0[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<3> DEC_X0[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<4> DEC_X0[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<5> DEC_X0[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<6> DEC_X0[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<7> DEC_X0[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<0> DEC_X1[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<1> DEC_X1[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<2> DEC_X1[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<3> DEC_X1[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<4> DEC_X1[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<5> DEC_X1[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<6> DEC_X1[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<7> DEC_X1[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    CNT_CORE_M8
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_CORE_M8 AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD 
+ PD_BUF PD_CVDDBUF PTSEL REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL 
+ VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] 
+ WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] 
+ XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] 
+ Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I PD:I PTSEL:I REDEN:I REDENB:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I 
*.PININFO XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I 
*.PININFO Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:O BIST2IO:O 
*.PININFO BLTRKWLDRV:O CKD:O DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O 
*.PININFO DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O DEC_X1[0]:O 
*.PININFO DEC_X1[1]:O DEC_X1[2]:O DEC_X1[3]:O DEC_X1[4]:O DEC_X1[5]:O 
*.PININFO DEC_X1[6]:O DEC_X1[7]:O DEC_X2[0]:O DEC_X2[1]:O DEC_X2[2]:O 
*.PININFO DEC_X2[3]:O DEC_X3[0]:O DEC_X3[1]:O DEC_X3[2]:O DEC_X3[3]:O 
*.PININFO DEC_X3[4]:O DEC_X3[5]:O DEC_X3[6]:O DEC_X3[7]:O DEC_Y[0]:O 
*.PININFO DEC_Y[1]:O DEC_Y[2]:O DEC_Y[3]:O DEC_Y[4]:O DEC_Y[5]:O DEC_Y[6]:O 
*.PININFO DEC_Y[7]:O PD_BUF:O PD_CVDDBUF:O RW_RE:O VHI:O VLO:O WLP_SAE:O 
*.PININFO WLP_SAEB:O YL[0]:O TK:B TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE_TK:B
MX0_PD<0> DEC_X0[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<1> DEC_X0[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<2> DEC_X0[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<3> DEC_X0[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<4> DEC_X0[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<5> DEC_X0[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<6> DEC_X0[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MX0_PD<7> DEC_X0[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<0> DEC_X1[0] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<1> DEC_X1[1] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<2> DEC_X1[2] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<3> DEC_X1[3] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<4> DEC_X1[4] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<5> DEC_X1[5] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<6> DEC_X1[6] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
MM0<7> DEC_X1[7] PD_BUF VSSI VSSI NCH L=60N W=400N M=1
XCDEC AX[0] AX[1] AX[2] AX[3] AX[4] AX[5] AX[6] AX[7] AX[8] AX[9] AX[10] 
+ BIST1B BIST2 CEB CEBM CK1B CK2 CKP CKPD CLK DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] EN ENC EN_DCLK PD REDEN REDENB RSC RW_RE 
+ VDDHD VDDI VSSI WEBXL WEBXL1B X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] 
+ X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] 
+ XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3] S1AHSF400W40_CDEC_M8M16
XCOTHERS AWT AWT2 BIST BIST1B BIST2 BIST2IO BLTRKWLDRV CK1B CK2 CKD CKP CKPD 
+ CLK EN ENC EN_DCLK PD PD_BUF PTSEL RSC RTSEL[0] RTSEL[1] TK TM TRKBL VDDHD 
+ VDDI VHI VLO VSSI WEB WEBM WEBXL WEBXL1B WLP_SAE WLP_SAEB WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2] S1AHSF400W40_COTH
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    CNT_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_CNT_SIM AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK CVDDHD CVDDI 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] 
+ FAD1[0] FAD1[1] FAD1[2] FAD1[3] FAD1[4] FAD1[5] FAD1[6] FAD1[7] FAD1[8] 
+ FAD1[9] FAD1[10] FAD2[0] FAD2[1] FAD2[2] FAD2[3] FAD2[4] FAD2[5] FAD2[6] 
+ FAD2[7] FAD2[8] FAD2[9] FAD2[10] HIT[0] HIT[1] PD PD_BUF PD_CVDDBUF PTSEL 
+ REDEN REDEN1 REDEN2 REDENB RSTB RTSEL[0] RTSEL[1] RW_RE SCLK SDIN SDOUT TK 
+ TM TRKBL VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAEB WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] 
+ X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] 
+ Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I CEB:I CEBM:I CLK:I FAD1[0]:I FAD1[1]:I FAD1[2]:I 
*.PININFO FAD1[3]:I FAD1[4]:I FAD1[5]:I FAD1[6]:I FAD1[7]:I FAD1[8]:I 
*.PININFO FAD1[9]:I FAD1[10]:I FAD2[0]:I FAD2[1]:I FAD2[2]:I FAD2[3]:I 
*.PININFO FAD2[4]:I FAD2[5]:I FAD2[6]:I FAD2[7]:I FAD2[8]:I FAD2[9]:I 
*.PININFO FAD2[10]:I PD:I PTSEL:I REDEN:I REDEN1:I REDEN2:I REDENB:I RSTB:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I SCLK:I SDIN:I TM:I WEB:I WEBM:I WTSEL[0]:I 
*.PININFO WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I 
*.PININFO X[6]:I X[7]:I X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I 
*.PININFO XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I 
*.PININFO Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I AWT2:B 
*.PININFO BIST2IO:B BLTRKWLDRV:B CKD:B CVDDHD:B CVDDI:B DEC_X0[0]:B 
*.PININFO DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B DEC_X0[5]:B 
*.PININFO DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B DEC_X1[2]:B 
*.PININFO DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B DEC_X1[7]:B 
*.PININFO DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B DEC_X3[0]:B 
*.PININFO DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B DEC_X3[4]:B DEC_X3[5]:B 
*.PININFO DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B 
*.PININFO DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B DEC_Y[7]:B HIT[0]:B HIT[1]:B 
*.PININFO PD_BUF:B PD_CVDDBUF:B RW_RE:B SDOUT:B TK:B TRKBL:B VDDHD:B VDDI:B 
*.PININFO VHI:B VLO:B VSSI:B WLP_SAE:B WLP_SAEB:B WLP_SAE_TK:B YL[0]:B
XI39 NET0539 NET0549 NET0160 NET0523 NET0384 NET0537 NET0495 NET0165 NET0517 
+ NET089[0] NET089[1] NET089[2] NET089[3] NET089[4] NET089[5] NET089[6] 
+ NET089[7] NET0518[0] NET0518[1] NET0518[2] NET0518[3] NET0518[4] NET0518[5] 
+ NET0518[6] NET0518[7] NET0572[0] NET0572[1] NET0572[2] NET0572[3] NET0192[0] 
+ NET0192[1] NET0192[2] NET0192[3] NET0192[4] NET0192[5] NET0192[6] NET0192[7] 
+ NET0531[0] NET0531[1] NET0531[2] NET0531[3] NET092[0] NET092[1] NET092[2] 
+ NET092[3] NET0157 NET0145 NET082 NET099 NET0133 NET093 NET0502[0] NET0502[1] 
+ NET0129 NET0127 NET0560 NET097 NET0570 NET098 NET0554 NET0190 NET0113 
+ NET0544 NET0540 NET0103 NET0199 NET0548 NET0526[0] NET0526[1] NET0526[2] 
+ NET0178[0] NET0178[1] NET0178[2] NET0178[3] NET0178[4] NET0178[5] NET0178[6] 
+ NET0178[7] NET0178[8] NET0178[9] NET0178[10] NET0507[0] NET0507[1] 
+ NET0507[2] NET0507[3] NET0507[4] NET0507[5] NET0507[6] NET0507[7] NET0507[8] 
+ NET0507[9] NET0507[10] NET0150[0] NET0150[1] NET0569 NET0186 NET0138 
+ NET0161[0] NET0161[1] NET070 NET0505 S1AHSF400W40_CNT_CORE_F_M16
XI40 NET0410 NET0387 NET0409 NET0128 NET0153 NET0408 NET0407 NET0115 NET0406 
+ NET0413[0] NET0413[1] NET0413[2] NET0413[3] NET0413[4] NET0413[5] NET0413[6] 
+ NET0413[7] NET0424[0] NET0424[1] NET0424[2] NET0424[3] NET0424[4] NET0424[5] 
+ NET0424[6] NET0424[7] NET0426[0] NET0426[1] NET0426[2] NET0426[3] NET0428[0] 
+ NET0428[1] NET0428[2] NET0428[3] NET0428[4] NET0428[5] NET0428[6] NET0428[7] 
+ NET0427[0] NET0427[1] NET0427[2] NET0427[3] NET0415[0] NET0415[1] NET0415[2] 
+ NET0415[3] NET0176 NET0423 NET0429 NET0425 NET0432 NET0198 NET0417[0] 
+ NET0417[1] NET0422 NET0416 NET0110 NET0414 NET0412 NET0411 NET0421 NET0420 
+ NET0393 NET096 NET0191 NET0419 NET0418 NET0124 NET0189[0] NET0189[1] 
+ NET0189[2] NET0182[0] NET0182[1] NET0182[2] NET0182[3] NET0182[4] NET0182[5] 
+ NET0182[6] NET0182[7] NET0182[8] NET0182[9] NET0182[10] NET0430[0] 
+ NET0430[1] NET0430[2] NET0430[3] NET0430[4] NET0430[5] NET0430[6] NET0430[7] 
+ NET0430[8] NET0430[9] NET0430[10] NET081[0] NET081[1] NET091 NET0397 NET0431 
+ NET0107[0] NET0107[1] NET0170 NET0177 S1AHSF400W40_CNT_CORE_F_M8
XI38 NET0453 NET0433 NET0452 NET0451 NET0458 NET0450 NET0448 NET0471 NET0447 
+ NET0474[0] NET0474[1] NET0474[2] NET0474[3] NET0474[4] NET0474[5] NET0474[6] 
+ NET0474[7] NET0476[0] NET0476[1] NET0476[2] NET0476[3] NET0476[4] NET0476[5] 
+ NET0476[6] NET0476[7] NET0477[0] NET0477[1] NET0477[2] NET0477[3] NET0478[0] 
+ NET0478[1] NET0478[2] NET0478[3] NET0478[4] NET0478[5] NET0478[6] NET0478[7] 
+ NET0475[0] NET0475[1] NET0475[2] NET0475[3] NET0470[0] NET0470[1] NET0470[2] 
+ NET0470[3] NET0446 NET0468 NET0469 NET0473 NET0449 NET0434 NET0462[0] 
+ NET0462[1] NET0467 NET0466 NET0445 NET0456 NET0455 NET0454 NET0465 NET0464 
+ NET0435 NET0444 NET0443 NET0463 NET0460 NET0461 NET0472[0] NET0472[1] 
+ NET0472[2] NET0442[0] NET0442[1] NET0442[2] NET0442[3] NET0442[4] NET0442[5] 
+ NET0442[6] NET0442[7] NET0442[8] NET0442[9] NET0442[10] NET0457[0] 
+ NET0457[1] NET0457[2] NET0457[3] NET0457[4] NET0457[5] NET0457[6] NET0457[7] 
+ NET0457[8] NET0457[9] NET0457[10] NET0441[0] NET0441[1] NET0440 NET0439 
+ NET0459 NET0438[0] NET0438[1] NET0437 NET0436 S1AHSF400W40_CNT_CORE_F_M4
XI35 NET0496 NET071 NET0149 NET0520 NET0141 NET079 NET0482 NET0200 NET0123 
+ NET0551[0] NET0551[1] NET0551[2] NET0551[3] NET0551[4] NET0551[5] NET0551[6] 
+ NET0551[7] NET073[0] NET073[1] NET073[2] NET073[3] NET073[4] NET073[5] 
+ NET073[6] NET073[7] NET0204[0] NET0204[1] NET0204[2] NET0204[3] NET0553[0] 
+ NET0553[1] NET0553[2] NET0553[3] NET0553[4] NET0553[5] NET0553[6] NET0553[7] 
+ NET0134[0] NET0134[1] NET0134[2] NET0134[3] NET0506[0] NET0506[1] NET0506[2] 
+ NET0506[3] NET0135 NET0126 NET0494 NET0562 NET0163 NET0203 NET090[0] 
+ NET090[1] NET0125 NET0575 NET0202 NET0132 NET085 NET0187 NET077 NET087 
+ NET0534 NET083 NET095 NET0512 NET0114 NET0513 NET0556[0] NET0556[1] 
+ NET0556[2] NET0195[0] NET0195[1] NET0195[2] NET0195[3] NET0195[4] NET0195[5] 
+ NET0195[6] NET0195[7] NET0195[8] NET0195[9] NET0195[10] NET0541[0] 
+ NET0541[1] NET0541[2] NET0541[3] NET0541[4] NET0541[5] NET0541[6] NET0541[7] 
+ NET0541[8] NET0541[9] NET0541[10] NET0117[0] NET0117[1] NET0532 NET078 
+ NET0183 NET0533[0] NET0533[1] NET0206 NET0205 S1AHSF400W40_CNT_CORE_F_M16_BIST
XI36 NET088 NET0159 NET069 NET0574 NET0555 NET0487 NET0535 NET0489 NET0571 
+ NET0558[0] NET0558[1] NET0558[2] NET0558[3] NET0558[4] NET0558[5] NET0558[6] 
+ NET0558[7] NET0168[0] NET0168[1] NET0168[2] NET0168[3] NET0168[4] NET0168[5] 
+ NET0168[6] NET0168[7] NET0545[0] NET0545[1] NET0545[2] NET0545[3] NET0201[0] 
+ NET0201[1] NET0201[2] NET0201[3] NET0201[4] NET0201[5] NET0201[6] NET0201[7] 
+ NET0516[0] NET0516[1] NET0516[2] NET0516[3] NET0563[0] NET0563[1] NET0563[2] 
+ NET0563[3] NET0175 NET0514 NET0143 NET0573 NET0501 NET0522 NET0180[0] 
+ NET0180[1] NET0152 NET0144 NET080 NET0504 NET0546 NET0142 NET0521 NET0119 
+ NET0171 NET0566 NET0481 NET076 NET0515 NET0536 NET0106[0] NET0106[1] 
+ NET0106[2] NET0547[0] NET0547[1] NET0547[2] NET0547[3] NET0547[4] NET0547[5] 
+ NET0547[6] NET0547[7] NET0547[8] NET0547[9] NET0547[10] NET0109[0] 
+ NET0109[1] NET0109[2] NET0109[3] NET0109[4] NET0109[5] NET0109[6] NET0109[7] 
+ NET0109[8] NET0109[9] NET0109[10] NET0139[0] NET0139[1] NET0488 NET0169 
+ NET0561 NET0162[0] NET0162[1] NET0172 NET0122 S1AHSF400W40_CNT_CORE_F_M8_BIST
XI37 NET0184 NET0491 NET0100 NET0527 NET0528 NET0565 NET094 NET0550 NET0185 
+ NET0130[0] NET0130[1] NET0130[2] NET0130[3] NET0130[4] NET0130[5] NET0130[6] 
+ NET0130[7] NET0497[0] NET0497[1] NET0497[2] NET0497[3] NET0497[4] NET0497[5] 
+ NET0497[6] NET0497[7] NET0131[0] NET0131[1] NET0131[2] NET0131[3] NET0196[0] 
+ NET0196[1] NET0196[2] NET0196[3] NET0196[4] NET0196[5] NET0196[6] NET0196[7] 
+ NET0111[0] NET0111[1] NET0111[2] NET0111[3] NET0483[0] NET0483[1] NET0483[2] 
+ NET0483[3] NET0567 NET0179 NET0116 NET0568 NET0140 NET0112 NET0559[0] 
+ NET0559[1] NET0104 NET0181 NET0136 NET0108 NET0155 NET0490 NET0156 NET0500 
+ NET0154 NET086 NET0519 NET0498 NET0146 NET084 NET0530[0] NET0530[1] 
+ NET0530[2] NET0173[0] NET0173[1] NET0173[2] NET0173[3] NET0173[4] NET0173[5] 
+ NET0173[6] NET0173[7] NET0173[8] NET0173[9] NET0173[10] NET0564[0] 
+ NET0564[1] NET0564[2] NET0564[3] NET0564[4] NET0564[5] NET0564[6] NET0564[7] 
+ NET0564[8] NET0564[9] NET0564[10] NET0137[0] NET0137[1] NET0529 NET0508 
+ NET0174 NET0158[0] NET0158[1] NET0509 NET0557 S1AHSF400W40_CNT_CORE_F_M4_BIST
XI0 NET0305 NET0333 NET0304 NET0332 NET0331 NET0303 NET0302 NET0330 NET0301 
+ NET0328[0] NET0328[1] NET0328[2] NET0328[3] NET0328[4] NET0328[5] NET0328[6] 
+ NET0328[7] NET0327[0] NET0327[1] NET0327[2] NET0327[3] NET0327[4] NET0327[5] 
+ NET0327[6] NET0327[7] NET0289[0] NET0289[1] NET0289[2] NET0289[3] NET0318[0] 
+ NET0318[1] NET0318[2] NET0318[3] NET0318[4] NET0318[5] NET0318[6] NET0318[7] 
+ NET0324[0] NET0324[1] NET0324[2] NET0324[3] NET0323[0] NET0323[1] NET0323[2] 
+ NET0323[3] NET0300 NET0319 NET0326 NET0325 NET0310 NET0288 NET0322[0] 
+ NET0322[1] NET0317 NET0329 NET0299 NET0309 NET0308 NET0307 NET0315 NET0314 
+ NET0306 NET0298 NET0297 NET0313 NET0312 NET0321 NET0320[0] NET0320[1] 
+ NET0320[2] NET0296[0] NET0296[1] NET0296[2] NET0296[3] NET0296[4] NET0296[5] 
+ NET0296[6] NET0296[7] NET0296[8] NET0296[9] NET0296[10] NET0316[0] 
+ NET0316[1] NET0316[2] NET0316[3] NET0316[4] NET0316[5] NET0316[6] NET0316[7] 
+ NET0316[8] NET0316[9] NET0316[10] NET0295[0] NET0295[1] NET0294 NET0293 
+ NET0311 NET0292[0] NET0292[1] NET0291 NET0290 S1AHSF400W40_CNT_CORE_M16_BIST
XI7 NET0357 NET0334 NET0356 NET0335 NET0336 NET0355 NET0354 NET0337 NET0353 
+ NET0360[0] NET0360[1] NET0360[2] NET0360[3] NET0360[4] NET0360[5] NET0360[6] 
+ NET0360[7] NET0371[0] NET0371[1] NET0371[2] NET0371[3] NET0371[4] NET0371[5] 
+ NET0371[6] NET0371[7] NET0373[0] NET0373[1] NET0373[2] NET0373[3] NET0375[0] 
+ NET0375[1] NET0375[2] NET0375[3] NET0375[4] NET0375[5] NET0375[6] NET0375[7] 
+ NET0374[0] NET0374[1] NET0374[2] NET0374[3] NET0362[0] NET0362[1] NET0362[2] 
+ NET0362[3] NET0352 NET0370 NET0376 NET0372 NET0379 NET0339 NET0364[0] 
+ NET0364[1] NET0369 NET0363 NET0351 NET0361 NET0359 NET0358 NET0368 NET0367 
+ NET0340 NET0350 NET0349 NET0366 NET0365 NET0338 NET0348[0] NET0348[1] 
+ NET0348[2] NET0347[0] NET0347[1] NET0347[2] NET0347[3] NET0347[4] NET0347[5] 
+ NET0347[6] NET0347[7] NET0347[8] NET0347[9] NET0347[10] NET0377[0] 
+ NET0377[1] NET0377[2] NET0377[3] NET0377[4] NET0377[5] NET0377[6] NET0377[7] 
+ NET0377[8] NET0377[9] NET0377[10] NET0346[0] NET0346[1] NET0345 NET0344 
+ NET0378 NET0343[0] NET0343[1] NET0342 NET0341 S1AHSF400W40_CNT_CORE_M8_BIST
XI8 NET0262 NET0242 NET0261 NET0260 NET0267 NET0259 NET0257 NET0280 NET0256 
+ NET0283[0] NET0283[1] NET0283[2] NET0283[3] NET0283[4] NET0283[5] NET0283[6] 
+ NET0283[7] NET0285[0] NET0285[1] NET0285[2] NET0285[3] NET0285[4] NET0285[5] 
+ NET0285[6] NET0285[7] NET0286[0] NET0286[1] NET0286[2] NET0286[3] NET0287[0] 
+ NET0287[1] NET0287[2] NET0287[3] NET0287[4] NET0287[5] NET0287[6] NET0287[7] 
+ NET0284[0] NET0284[1] NET0284[2] NET0284[3] NET0279[0] NET0279[1] NET0279[2] 
+ NET0279[3] NET0255 NET0277 NET0278 NET0282 NET0258 NET0243 NET0271[0] 
+ NET0271[1] NET0276 NET0275 NET0254 NET0265 NET0264 NET0263 NET0274 NET0273 
+ NET0244 NET0253 NET0252 NET0272 NET0269 NET0270 NET0281[0] NET0281[1] 
+ NET0281[2] NET0251[0] NET0251[1] NET0251[2] NET0251[3] NET0251[4] NET0251[5] 
+ NET0251[6] NET0251[7] NET0251[8] NET0251[9] NET0251[10] NET0266[0] 
+ NET0266[1] NET0266[2] NET0266[3] NET0266[4] NET0266[5] NET0266[6] NET0266[7] 
+ NET0266[8] NET0266[9] NET0266[10] NET0250[0] NET0250[1] NET0249 NET0248 
+ NET0268 NET0247[0] NET0247[1] NET0246 NET0245 S1AHSF400W40_CNT_CORE_M4_BIST
XI34 NET029 NET064 NET0401 NET0395 NET068 NET0121 NET019 NET057 NET0118 
+ NET0403[0] NET0403[1] NET0403[2] NET0403[3] NET0403[4] NET0403[5] NET0403[6] 
+ NET0403[7] NET0147[0] NET0147[1] NET0147[2] NET0147[3] NET0147[4] NET0147[5] 
+ NET0147[6] NET0147[7] NET0148[0] NET0148[1] NET0148[2] NET0148[3] NET0404[0] 
+ NET0404[1] NET0404[2] NET0404[3] NET0404[4] NET0404[5] NET0404[6] NET0404[7] 
+ NET037[0] NET037[1] NET037[2] NET037[3] NET0396[0] NET0396[1] NET0396[2] 
+ NET0396[3] NET028 NET0405 NET036 NET025 NET0120 NET0105 NET032[0] NET032[1] 
+ NET054 NET059 NET053 NET018 NET0388 NET024 NET035 NET013 NET075 NET039 NET07 
+ NET0389 NET010 NET0398 NET030[0] NET030[1] NET030[2] NET056[0] NET056[1] 
+ NET056[2] NET056[3] NET056[4] NET056[5] NET056[6] NET056[7] NET056[8] 
+ NET056[9] NET056[10] NET050[0] NET050[1] NET050[2] NET050[3] NET050[4] 
+ NET050[5] NET050[6] NET050[7] NET050[8] NET050[9] NET050[10] NET042[0] 
+ NET042[1] NET065 NET038 NET058 NET044[0] NET044[1] NET063 NET020 
+ S1AHSF400W40_CNT_CORE_M4
XI33 NET0167 NET060 NET0166 NET0194 NET0193 NET022 NET0164 NET055 NET034 
+ NET0385[0] NET0385[1] NET0385[2] NET0385[3] NET0385[4] NET0385[5] NET0385[6] 
+ NET0385[7] NET046[0] NET046[1] NET046[2] NET046[3] NET046[4] NET046[5] 
+ NET046[6] NET046[7] NET0151[0] NET0151[1] NET0151[2] NET0151[3] NET031[0] 
+ NET031[1] NET031[2] NET031[3] NET031[4] NET031[5] NET031[6] NET031[7] 
+ NET021[0] NET021[1] NET021[2] NET021[3] NET0394[0] NET0394[1] NET0394[2] 
+ NET0394[3] NET048 NET041 NET0188 NET0386 NET011 NET0380 NET045[0] NET045[1] 
+ NET066 NET0383 NET051 NET043 NET0400 NET0381 NET017 NET052 NET015 NET0392 
+ NET072 NET033 NET0390 NET067 NET0101[0] NET0101[1] NET0101[2] NET0102[0] 
+ NET0102[1] NET0102[2] NET0102[3] NET0102[4] NET0102[5] NET0102[6] NET0102[7] 
+ NET0102[8] NET0102[9] NET0102[10] NET09[0] NET09[1] NET09[2] NET09[3] 
+ NET09[4] NET09[5] NET09[6] NET09[7] NET09[8] NET09[9] NET09[10] NET027[0] 
+ NET027[1] NET014 NET08 NET023 NET0382[0] NET0382[1] NET0399 NET0402 
+ S1AHSF400W40_CNT_CORE_M16
XI32 NET0219 NET062 NET0218 NET0197 NET026 NET0217 NET0216 NET0391 NET0215 
+ NET0222[0] NET0222[1] NET0222[2] NET0222[3] NET0222[4] NET0222[5] NET0222[6] 
+ NET0222[7] NET0233[0] NET0233[1] NET0233[2] NET0233[3] NET0233[4] NET0233[5] 
+ NET0233[6] NET0233[7] NET0235[0] NET0235[1] NET0235[2] NET0235[3] NET0237[0] 
+ NET0237[1] NET0237[2] NET0237[3] NET0237[4] NET0237[5] NET0237[6] NET0237[7] 
+ NET0236[0] NET0236[1] NET0236[2] NET0236[3] NET0224[0] NET0224[1] NET0224[2] 
+ NET0224[3] NET0214 NET0232 NET0238 NET0234 NET0241 NET040 NET0226[0] 
+ NET0226[1] NET0231 NET0225 NET0213 NET0223 NET0221 NET0220 NET0230 NET0229 
+ NET016 NET0212 NET0211 NET0228 NET0227 NET061 NET0210[0] NET0210[1] 
+ NET0210[2] NET0209[0] NET0209[1] NET0209[2] NET0209[3] NET0209[4] NET0209[5] 
+ NET0209[6] NET0209[7] NET0209[8] NET0209[9] NET0209[10] NET0239[0] 
+ NET0239[1] NET0239[2] NET0239[3] NET0239[4] NET0239[5] NET0239[6] NET0239[7] 
+ NET0239[8] NET0239[9] NET0239[10] NET0208[0] NET0208[1] NET0207 NET012 
+ NET0240 NET049[0] NET049[1] NET047 NET074 S1AHSF400W40_CNT_CORE_M8
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    DOUT
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_DOUT AWT AWTD GBL GBLB PD Q VDDHD VSSI WLP_SAEB
*.PININFO AWT:I AWTD:I PD:I WLP_SAEB:I Q:O GBL:B GBLB:B VDDHD:B VSSI:B
MP11 NET083 NET065 VDDHD VDDHD PCH L=60N W=1U M=3
MP0 GBLB GBL VDDHD VDDHD PCH L=60N W=360.0N M=1
MP6 VDDHD GBLB GBL VDDHD PCH L=60N W=360.0N M=1
MP7 VDDHD DLRSB GBLB VDDHD PCH L=60N W=1U M=6
MP8 GBL DLRSB VDDHD VDDHD PCH L=60N W=1U M=6
MP4 QBB QB VDDHD VDDHD PCH L=60N W=1.25U M=2
MP9 NET095 QBB VDDHD VDDHD PCH L=60N W=1.25U M=2
MP5 NET095 GBL VDDHD VDDHD PCH L=60N W=1.25U M=2
MP15 QBB GBLB VDDHD VDDHD PCH L=60N W=1.25U M=2
MP2 NET095 AWT QB VDDHD PCH L=60N W=1.25U M=4
MM0 QB AWT1B NET083 VDDHD PCH L=60N W=1U M=3
MN6 NET0127 NET065 VSSI VSSI NCH L=60N W=500N M=3
MN20 Z3 GBL Z2 VSSI NCH L=60N W=1.25U M=3
MM1 QB AWT NET0127 VSSI NCH L=60N W=500N M=3
MN8 Z2 AWT1B VSSI VSSI NCH L=60N W=1.25U M=3
MN21 QBB GBLB Z1 VSSI NCH L=60N W=1.25U M=2
MN22 Z1 QB VSSI VSSI NCH L=60N W=1.25U M=2
MN18 QB QBB Z3 VSSI NCH L=60N W=1.25U M=3
XI154 AWTD VSSI VDDHD AWTD1B S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.5U 
+ LP=0.06U M=1
XI153 AWTD1B VSSI VDDHD NET065 S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U 
+ LP=0.06U M=1
XI109 QB VSSI VDDHD Q S1AHSF400W40_AINV FN=4 WN=0.5U LN=0.06U FP=4 WP=1U LP=0.06U M=1
XINV3 WLP_SAEB VSSI VDDHD DLRSB S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U 
+ LP=0.06U M=1
XINV1 AWT VSSI VDDHD AWT1B S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    DIN
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_DIN AWTD BIST BWEB BWEBM CKD D DM GW GWB VDDHD VDDI VSSI
*.PININFO BIST:I BWEB:I BWEBM:I CKD:I D:I DM:I AWTD:O GW:O GWB:O VDDHD:B 
*.PININFO VDDI:B VSSI:B
XI324 CKD1B VSSI VSSI VDDHD VDDHD CKD2 S1AHSF400W40_INV_BULK FN=1 WN=0.6U LN=0.06U FP=1 
+ WP=1.2U LP=0.06U M=1
XI323 CKD VSSI VSSI VDDHD VDDHD CKD1B S1AHSF400W40_INV_BULK FN=1 WN=0.4U LN=0.06U FP=1 
+ WP=0.8U LP=0.06U M=1
XI326 BIST1B VSSI VSSI VDDHD VDDHD BIST2 S1AHSF400W40_INV_BULK FN=1 WN=0.6U LN=0.06U FP=1 
+ WP=1.2U LP=0.06U M=1
XI325 BIST VSSI VSSI VDDHD VDDHD BIST1B S1AHSF400W40_INV_BULK FN=1 WN=0.4U LN=0.06U FP=1 
+ WP=0.8U LP=0.06U M=1
MM51 DXL3B_AND DXL2 VDDHD VDDHD PCH L=60N W=500N M=2
MM52 DXL2_AND DXL1B VDDHD VDDHD PCH L=60N W=500N M=2
MM53 DXL2_AND BXL1B VDDHD VDDHD PCH L=60N W=500N M=2
MM54 DXL3B_AND BXL1B VDDHD VDDHD PCH L=60N W=500N M=2
MM26 VDDHD CKD2 Z9 VDDHD PCH L=120.0N W=600N M=1
MM38 VDDHD CKD2 Z13 VDDHD PCH L=120.0N W=600N M=1
MM39 VDDHD BXL1B Z16 VDDHD PCH L=120.0N W=600N M=1
MM40 BXL CKD1B Z16 VDDHD PCH L=120.0N W=600N M=1
MM22 Z21 D VDDHD VDDHD PCH L=120.0N W=600N M=1
MM27 DXL DXB Z9 VDDHD PCH L=120.0N W=600N M=1
MM29 DXL CKD1B Z6 VDDHD PCH L=120.0N W=600N M=1
MM24 D_BIST BIST1B Z22 VDDHD PCH L=120.0N W=600N M=1
MM23 D_BIST BIST2 Z21 VDDHD PCH L=120.0N W=600N M=1
MM41 BXL BXB Z13 VDDHD PCH L=120.0N W=600N M=1
MP2 AWTD DX Z18 VDDHD PCH L=60N W=800N M=1
MP3 Z18 BXB VDDHD VDDHD PCH L=60N W=800N M=1
MP18 Z25 BWEB VDDHD VDDHD PCH L=120.0N W=600N M=1
MP19 B_BIST BIST2 Z25 VDDHD PCH L=120.0N W=600N M=1
MP4 Z19 BX VDDHD VDDHD PCH L=60N W=800N M=1
MP5 AWTD DXB Z19 VDDHD PCH L=60N W=800N M=1
MP16 B_BIST BIST1B Z26 VDDHD PCH L=120.0N W=600N M=1
MM28 VDDHD DXL1B Z6 VDDHD PCH L=120.0N W=600N M=1
MM25 Z22 DM VDDHD VDDHD PCH L=120.0N W=600N M=1
MP25 Z26 BWEBM VDDHD VDDHD PCH L=120.0N W=600N M=1
MP10 DXL2_AND CKD2 VDDHD VDDHD PCH L=60N W=500N M=2
MP1 DXL3B_AND CKD2 VDDHD VDDHD PCH L=60N W=500N M=2
MM35 DXL CKD2 Z7 VSSI NCH L=120.0N W=300N M=1
MN33 DXL3B_AND DXL2 Z2 VSSI NCH L=60N W=2U M=1
MM33 D_BIST BIST2 Z24 VSSI NCH L=120.0N W=300N M=1
MM32 Z24 DM VSSI VSSI NCH L=120.0N W=300N M=1
MM36 VSSI CKD1B Z11 VSSI NCH L=120.0N W=300N M=1
MM34 DXL DXB Z11 VSSI NCH L=120.0N W=300N M=1
MM31 Z23 D VSSI VSSI NCH L=120.0N W=300N M=1
MM30 D_BIST BIST1B Z23 VSSI NCH L=120.0N W=300N M=1
MN2 Z2 CKD2 Z1 VSSI NCH L=60N W=1U M=4
MN27 B_BIST BIST2 Z28 VSSI NCH L=120.0N W=300N M=1
MM37 VSSI DXL1B Z7 VSSI NCH L=120.0N W=300N M=1
MM43 VSSI CKD1B Z15 VSSI NCH L=120.0N W=300N M=1
MM42 BXL BXB Z15 VSSI NCH L=120.0N W=300N M=1
MN13 Z20 DXB VSSI VSSI NCH L=60N W=400N M=1
MN6 AWTD DX Z20 VSSI NCH L=60N W=400N M=1
MN16 Z28 BWEBM VSSI VSSI NCH L=120.0N W=300N M=1
MN5 AWTD BXB Z20 VSSI NCH L=60N W=400N M=1
MN4 Z20 BX VSSI VSSI NCH L=60N W=400N M=1
MM44 VSSI BXL1B Z14 VSSI NCH L=120.0N W=300N M=1
MM45 BXL CKD2 Z14 VSSI NCH L=120.0N W=300N M=1
MN19 B_BIST BIST1B Z27 VSSI NCH L=120.0N W=300N M=1
MN7 Z1 BXL1B VSSI VSSI NCH L=60N W=1U M=6
MN17 Z27 BWEB VSSI VSSI NCH L=120.0N W=300N M=1
MN1 DXL2_AND DXL1B Z2 VSSI NCH L=60N W=1U M=2
XINV00 D_BIST VSSI VDDHD DX S1AHSF400W40_AINV FN=1 WN=0.3U LN=120N FP=1 WP=0.3U LP=120N 
+ M=1
XINV05 DXL1B VSSI VDDHD DXL2 S1AHSF400W40_AINV FN=2 WN=0.3U LN=0.06U FP=2 WP=0.6U 
+ LP=0.06U M=1
XINV07 DXL3B_AND VSSI VDDHD GW S1AHSF400W40_AINV FN=6 WN=0.8U LN=0.06U FP=6 WP=1.6U 
+ LP=0.06U M=1
XI317 DXL2_AND VSSI VDDHD GWB S1AHSF400W40_AINV FN=6 WN=0.8U LN=0.06U FP=6 WP=1.6U 
+ LP=0.06U M=1
XI319 BXL VSSI VDDHD BXL1B S1AHSF400W40_AINV FN=2 WN=0.3U LN=0.06U FP=2 WP=0.6U LP=0.06U 
+ M=1
XI315 B_BIST VSSI VDDHD BX S1AHSF400W40_AINV FN=1 WN=0.3U LN=120N FP=1 WP=0.3U LP=120N M=1
XI318 DXL VSSI VDDHD DXL1B S1AHSF400W40_AINV FN=2 WN=0.3U LN=0.06U FP=2 WP=0.6U LP=0.06U 
+ M=1
XINV01 DX VSSI VDDHD DXB S1AHSF400W40_AINV FN=1 WN=0.3U LN=120N FP=1 WP=0.3U LP=120N M=1
XI316 BX VSSI VDDHD BXB S1AHSF400W40_AINV FN=1 WN=0.3U LN=120N FP=1 WP=0.3U LP=120N M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    IO
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_IO AWT BIST BWEB BWEBM CKD D DM GBL GBLB GW GWB PD Q VDDHD VDDI VSSI 
+ WLP_SAEB
*.PININFO AWT:I BIST:I BWEB:I BWEBM:I CKD:I D:I DM:I PD:I WLP_SAEB:I GW:O 
*.PININFO GWB:O Q:O GBL:B GBLB:B VDDHD:B VDDI:B VSSI:B
XDOUT AWT AWTD GBL GBLB PD Q VDDHD VSSI WLP_SAEB S1AHSF400W40_DOUT
XDIN AWTD BIST BWEB BWEBM CKD D DM GW GWB VDDHD VDDI VSSI S1AHSF400W40_DIN
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    IO_M16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_IO_M16 AWT2 BIST2IO BWEB BWEBM CKD D DM GBL GBLB GW GWB PD_BUF Q VDDHD 
+ VDDI VSSI WLP_SAEB
*.PININFO AWT2:I BIST2IO:I BWEB:I BWEBM:I CKD:I D:I DM:I PD_BUF:I WLP_SAEB:I 
*.PININFO GW:O GWB:O Q:O GBL:B GBLB:B VDDHD:B VDDI:B VSSI:B
MN7 Q PD_BUF VSSI VSSI NCH L=60N W=500N M=1
XIO AWT2 BIST2IO BWEB BWEBM CKD D DM GBL GBLB GW GWB PD_BUF Q VDDHD VDDI VSSI 
+ WLP_SAEB S1AHSF400W40_IO
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    IO_M8
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_IO_M8 AWT2 BIST2IO BWEB BWEBM CKD D DM GBL GBLB GW GWB PD_BUF Q VDDHD 
+ VDDI VSSI WLP_SAEB
*.PININFO AWT2:I BIST2IO:I BWEB:I BWEBM:I CKD:I D:I DM:I PD_BUF:I WLP_SAEB:I 
*.PININFO GW:O GWB:O Q:O GBL:B GBLB:B VDDHD:B VDDI:B VSSI:B
MN7 Q PD_BUF VSSI VSSI NCH L=60N W=500N M=1
XIO AWT2 BIST2IO BWEB BWEBM CKD D DM GBL GBLB GW GWB PD_BUF Q VDDHD VDDI VSSI 
+ WLP_SAEB S1AHSF400W40_IO
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    IO_M4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_IO_M4 AWT2 BIST2IO BWEB BWEBM CKD D DM GBL GBLB GW GWB PD_BUF Q VDDHD 
+ VDDI VSSI WLP_SAEB
*.PININFO AWT2:I BIST2IO:I BWEB:I BWEBM:I CKD:I D:I DM:I PD_BUF:I WLP_SAEB:I 
*.PININFO GW:O GWB:O Q:O GBL:B GBLB:B VDDHD:B VDDI:B VSSI:B
MN7 Q PD_BUF VSSI VSSI NCH L=60N W=500N M=1
XIO AWT2 BIST2IO BWEB BWEBM CKD D DM GBL GBLB GW GWB PD_BUF Q VDDHD VDDI VSSI 
+ WLP_SAEB S1AHSF400W40_IO
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    IO_LD_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_IO_LD_SIM AWT2_LT AWT2_RT BIST2IO_LT BIST2IO_RT CKD_LT CKD_RT 
+ PD_BUF_LT PD_BUF_RT VDDHD VDDI VSSI WLP_SAEB_LT WLP_SAEB_RT
*.PININFO AWT2_LT:B AWT2_RT:B BIST2IO_LT:B BIST2IO_RT:B CKD_LT:B CKD_RT:B 
*.PININFO PD_BUF_LT:B PD_BUF_RT:B VDDHD:B VDDI:B VSSI:B WLP_SAEB_LT:B 
*.PININFO WLP_SAEB_RT:B
XIO_M16 NET03 NET01 NET011 NET06 NET010 NET09 NET012 NET07 NET04 NET013 NET027 
+ NET05 NET02 NET030 NET028 NET029 NET08 S1AHSF400W40_IO_M16
XIO_M8 NET035 NET034 NET039 NET038 NET031 NET037 NET036 NET033 NET042 NET040 
+ NET044 NET032 NET041 NET047 NET045 NET046 NET043 S1AHSF400W40_IO_M8
XIO_M4 NET052 NET051 NET056 NET055 NET048 NET054 NET053 NET050 NET059 NET057 
+ NET061 NET049 NET058 NET064 NET062 NET063 NET060 S1AHSF400W40_IO_M4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    IO_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_IO_SIM AWT2_LT AWT2_RT BIST2IO_LT BIST2IO_RT BWEBM_BT BWEB_BT CKD_LT 
+ CKD_RT DM_BT D_BT GBLB_TP GBL_TP GWB_TP GW_TP PD_BUF_LT PD_BUF_RT Q_BT VDDHD 
+ VDDI VSSI WLP_SAEB_LT WLP_SAEB_RT
*.PININFO AWT2_LT:B AWT2_RT:B BIST2IO_LT:B BIST2IO_RT:B BWEBM_BT:B BWEB_BT:B 
*.PININFO CKD_LT:B CKD_RT:B DM_BT:B D_BT:B GBLB_TP:B GBL_TP:B GWB_TP:B GW_TP:B 
*.PININFO PD_BUF_LT:B PD_BUF_RT:B Q_BT:B VDDHD:B VDDI:B VSSI:B WLP_SAEB_LT:B 
*.PININFO WLP_SAEB_RT:B
XIO_M16 NET062 NET013 NET066 NET065 NET012 NET064 NET063 NET018 NET069 NET067 
+ NET071 NET02 NET068 NET074 NET072 NET073 NET070 S1AHSF400W40_IO_M16
XIO_M8 NET079 NET078 NET083 NET082 NET075 NET081 NET080 NET077 NET086 NET084 
+ NET088 NET076 NET085 NET091 NET089 NET090 NET087 S1AHSF400W40_IO_M8
XIO_M4 NET096 NET095 NET0100 NET099 NET092 NET06 NET020 NET094 NET0103 NET023 
+ NET022 NET093 NET0102 NET016 NET019 NET0107 NET017 S1AHSF400W40_IO_M4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MCB_2X4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_2X4 BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB 
+ GW GWB VDDI VSSI WL[0] WL[1]
*.PININFO WL[0]:I WL[1]:I BL[0]:B BL[1]:B BL[2]:B BL[3]:B BLB[0]:B BLB[1]:B 
*.PININFO BLB[2]:B BLB[3]:B GBL:B GBLB:B GW:B GWB:B VDDI:B VSSI:B
XMCB_0<0> BL[0] BLB[0] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<1> BL[1] BLB[1] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<2> BL[2] BLB[2] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<3> BL[3] BLB[3] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_1<0> BL[0] BLB[0] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<1> BL[1] BLB[1] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<2> BL[2] BLB[2] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<3> BL[3] BLB[3] VDDI VSSI WL[1] S1AHSF400W40_MCB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    MCB_32X4_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_32X4_CHAR BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL 
+ GBLB GW GWB VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] 
+ WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] 
+ WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] 
+ WL[31]
*.PININFO WL[0]:I WL[1]:I WL[2]:I WL[3]:I WL[4]:I WL[5]:I WL[6]:I WL[7]:I 
*.PININFO WL[8]:I WL[9]:I WL[10]:I WL[11]:I WL[12]:I WL[13]:I WL[14]:I 
*.PININFO WL[15]:I WL[16]:I WL[17]:I WL[18]:I WL[19]:I WL[20]:I WL[21]:I 
*.PININFO WL[22]:I WL[23]:I WL[24]:I WL[25]:I WL[26]:I WL[27]:I WL[28]:I 
*.PININFO WL[29]:I WL[30]:I WL[31]:I BL[0]:B BL[1]:B BL[2]:B BL[3]:B BLB[0]:B 
*.PININFO BLB[1]:B BLB[2]:B BLB[3]:B GBL:B GBLB:B GW:B GWB:B VDDI:B VSSI:B
XMCB_2X4<0> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_2X4<1> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[2] WL[3] S1AHSF400W40_MCB_2X4
XMCB_2X4<2> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[4] WL[5] S1AHSF400W40_MCB_2X4
XMCB_2X4<3> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[6] WL[7] S1AHSF400W40_MCB_2X4
XMCB_2X4<4> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[8] WL[9] S1AHSF400W40_MCB_2X4
XMCB_2X4<5> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[10] WL[11] S1AHSF400W40_MCB_2X4
XMCB_2X4<6> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[12] WL[13] S1AHSF400W40_MCB_2X4
XMCB_2X4<7> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[14] WL[15] S1AHSF400W40_MCB_2X4
XMCB_2X4<8> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[16] WL[17] S1AHSF400W40_MCB_2X4
XMCB_2X4<9> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[18] WL[19] S1AHSF400W40_MCB_2X4
XMCB_2X4<10> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[20] WL[21] S1AHSF400W40_MCB_2X4
XMCB_2X4<11> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[22] WL[23] S1AHSF400W40_MCB_2X4
XMCB_2X4<12> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[24] WL[25] S1AHSF400W40_MCB_2X4
XMCB_2X4<13> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[26] WL[27] S1AHSF400W40_MCB_2X4
XMCB_2X4<14> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[28] WL[29] S1AHSF400W40_MCB_2X4
XMCB_2X4<15> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[30] WL[31] S1AHSF400W40_MCB_2X4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    MCB_64X4_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_64X4_CHAR BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL 
+ GBLB GW GWB VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] 
+ WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] 
+ WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] 
+ WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] 
+ WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] 
+ WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63]
*.PININFO WL[0]:I WL[1]:I WL[2]:I WL[3]:I WL[4]:I WL[5]:I WL[6]:I WL[7]:I 
*.PININFO WL[8]:I WL[9]:I WL[10]:I WL[11]:I WL[12]:I WL[13]:I WL[14]:I 
*.PININFO WL[15]:I WL[16]:I WL[17]:I WL[18]:I WL[19]:I WL[20]:I WL[21]:I 
*.PININFO WL[22]:I WL[23]:I WL[24]:I WL[25]:I WL[26]:I WL[27]:I WL[28]:I 
*.PININFO WL[29]:I WL[30]:I WL[31]:I WL[32]:I WL[33]:I WL[34]:I WL[35]:I 
*.PININFO WL[36]:I WL[37]:I WL[38]:I WL[39]:I WL[40]:I WL[41]:I WL[42]:I 
*.PININFO WL[43]:I WL[44]:I WL[45]:I WL[46]:I WL[47]:I WL[48]:I WL[49]:I 
*.PININFO WL[50]:I WL[51]:I WL[52]:I WL[53]:I WL[54]:I WL[55]:I WL[56]:I 
*.PININFO WL[57]:I WL[58]:I WL[59]:I WL[60]:I WL[61]:I WL[62]:I WL[63]:I 
*.PININFO BL[0]:B BL[1]:B BL[2]:B BL[3]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B 
*.PININFO GBL:B GBLB:B GW:B GWB:B VDDI:B VSSI:B
XMCB_2X4<0> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_2X4<1> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[2] WL[3] S1AHSF400W40_MCB_2X4
XMCB_2X4<2> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[4] WL[5] S1AHSF400W40_MCB_2X4
XMCB_2X4<3> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[6] WL[7] S1AHSF400W40_MCB_2X4
XMCB_2X4<4> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[8] WL[9] S1AHSF400W40_MCB_2X4
XMCB_2X4<5> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[10] WL[11] S1AHSF400W40_MCB_2X4
XMCB_2X4<6> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[12] WL[13] S1AHSF400W40_MCB_2X4
XMCB_2X4<7> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[14] WL[15] S1AHSF400W40_MCB_2X4
XMCB_2X4<8> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[16] WL[17] S1AHSF400W40_MCB_2X4
XMCB_2X4<9> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[18] WL[19] S1AHSF400W40_MCB_2X4
XMCB_2X4<10> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[20] WL[21] S1AHSF400W40_MCB_2X4
XMCB_2X4<11> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[22] WL[23] S1AHSF400W40_MCB_2X4
XMCB_2X4<12> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[24] WL[25] S1AHSF400W40_MCB_2X4
XMCB_2X4<13> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[26] WL[27] S1AHSF400W40_MCB_2X4
XMCB_2X4<14> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[28] WL[29] S1AHSF400W40_MCB_2X4
XMCB_2X4<15> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[30] WL[31] S1AHSF400W40_MCB_2X4
XMCB_2X4<16> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[32] WL[33] S1AHSF400W40_MCB_2X4
XMCB_2X4<17> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[34] WL[35] S1AHSF400W40_MCB_2X4
XMCB_2X4<18> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[36] WL[37] S1AHSF400W40_MCB_2X4
XMCB_2X4<19> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[38] WL[39] S1AHSF400W40_MCB_2X4
XMCB_2X4<20> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[40] WL[41] S1AHSF400W40_MCB_2X4
XMCB_2X4<21> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[42] WL[43] S1AHSF400W40_MCB_2X4
XMCB_2X4<22> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[44] WL[45] S1AHSF400W40_MCB_2X4
XMCB_2X4<23> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[46] WL[47] S1AHSF400W40_MCB_2X4
XMCB_2X4<24> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[48] WL[49] S1AHSF400W40_MCB_2X4
XMCB_2X4<25> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[50] WL[51] S1AHSF400W40_MCB_2X4
XMCB_2X4<26> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[52] WL[53] S1AHSF400W40_MCB_2X4
XMCB_2X4<27> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[54] WL[55] S1AHSF400W40_MCB_2X4
XMCB_2X4<28> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[56] WL[57] S1AHSF400W40_MCB_2X4
XMCB_2X4<29> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[58] WL[59] S1AHSF400W40_MCB_2X4
XMCB_2X4<30> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[60] WL[61] S1AHSF400W40_MCB_2X4
XMCB_2X4<31> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[62] WL[63] S1AHSF400W40_MCB_2X4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    MCB_128X4_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_128X4_CHAR BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL 
+ GBLB GW GWB VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] 
+ WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] 
+ WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] 
+ WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] 
+ WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] 
+ WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] 
+ WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] WL[72] WL[73] WL[74] 
+ WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] WL[83] WL[84] WL[85] 
+ WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] WL[94] WL[95] WL[96] 
+ WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] WL[104] WL[105] WL[106] 
+ WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] WL[113] WL[114] WL[115] 
+ WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] WL[122] WL[123] WL[124] 
+ WL[125] WL[126] WL[127]
*.PININFO WL[0]:I WL[1]:I WL[2]:I WL[3]:I WL[4]:I WL[5]:I WL[6]:I WL[7]:I 
*.PININFO WL[8]:I WL[9]:I WL[10]:I WL[11]:I WL[12]:I WL[13]:I WL[14]:I 
*.PININFO WL[15]:I WL[16]:I WL[17]:I WL[18]:I WL[19]:I WL[20]:I WL[21]:I 
*.PININFO WL[22]:I WL[23]:I WL[24]:I WL[25]:I WL[26]:I WL[27]:I WL[28]:I 
*.PININFO WL[29]:I WL[30]:I WL[31]:I WL[32]:I WL[33]:I WL[34]:I WL[35]:I 
*.PININFO WL[36]:I WL[37]:I WL[38]:I WL[39]:I WL[40]:I WL[41]:I WL[42]:I 
*.PININFO WL[43]:I WL[44]:I WL[45]:I WL[46]:I WL[47]:I WL[48]:I WL[49]:I 
*.PININFO WL[50]:I WL[51]:I WL[52]:I WL[53]:I WL[54]:I WL[55]:I WL[56]:I 
*.PININFO WL[57]:I WL[58]:I WL[59]:I WL[60]:I WL[61]:I WL[62]:I WL[63]:I 
*.PININFO WL[64]:I WL[65]:I WL[66]:I WL[67]:I WL[68]:I WL[69]:I WL[70]:I 
*.PININFO WL[71]:I WL[72]:I WL[73]:I WL[74]:I WL[75]:I WL[76]:I WL[77]:I 
*.PININFO WL[78]:I WL[79]:I WL[80]:I WL[81]:I WL[82]:I WL[83]:I WL[84]:I 
*.PININFO WL[85]:I WL[86]:I WL[87]:I WL[88]:I WL[89]:I WL[90]:I WL[91]:I 
*.PININFO WL[92]:I WL[93]:I WL[94]:I WL[95]:I WL[96]:I WL[97]:I WL[98]:I 
*.PININFO WL[99]:I WL[100]:I WL[101]:I WL[102]:I WL[103]:I WL[104]:I WL[105]:I 
*.PININFO WL[106]:I WL[107]:I WL[108]:I WL[109]:I WL[110]:I WL[111]:I 
*.PININFO WL[112]:I WL[113]:I WL[114]:I WL[115]:I WL[116]:I WL[117]:I 
*.PININFO WL[118]:I WL[119]:I WL[120]:I WL[121]:I WL[122]:I WL[123]:I 
*.PININFO WL[124]:I WL[125]:I WL[126]:I WL[127]:I BL[0]:B BL[1]:B BL[2]:B 
*.PININFO BL[3]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B GBL:B GBLB:B GW:B GWB:B 
*.PININFO VDDI:B VSSI:B
XMCB_2X4<0> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_2X4<1> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[2] WL[3] S1AHSF400W40_MCB_2X4
XMCB_2X4<2> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[4] WL[5] S1AHSF400W40_MCB_2X4
XMCB_2X4<3> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[6] WL[7] S1AHSF400W40_MCB_2X4
XMCB_2X4<4> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[8] WL[9] S1AHSF400W40_MCB_2X4
XMCB_2X4<5> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[10] WL[11] S1AHSF400W40_MCB_2X4
XMCB_2X4<6> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[12] WL[13] S1AHSF400W40_MCB_2X4
XMCB_2X4<7> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[14] WL[15] S1AHSF400W40_MCB_2X4
XMCB_2X4<8> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[16] WL[17] S1AHSF400W40_MCB_2X4
XMCB_2X4<9> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[18] WL[19] S1AHSF400W40_MCB_2X4
XMCB_2X4<10> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[20] WL[21] S1AHSF400W40_MCB_2X4
XMCB_2X4<11> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[22] WL[23] S1AHSF400W40_MCB_2X4
XMCB_2X4<12> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[24] WL[25] S1AHSF400W40_MCB_2X4
XMCB_2X4<13> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[26] WL[27] S1AHSF400W40_MCB_2X4
XMCB_2X4<14> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[28] WL[29] S1AHSF400W40_MCB_2X4
XMCB_2X4<15> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[30] WL[31] S1AHSF400W40_MCB_2X4
XMCB_2X4<16> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[32] WL[33] S1AHSF400W40_MCB_2X4
XMCB_2X4<17> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[34] WL[35] S1AHSF400W40_MCB_2X4
XMCB_2X4<18> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[36] WL[37] S1AHSF400W40_MCB_2X4
XMCB_2X4<19> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[38] WL[39] S1AHSF400W40_MCB_2X4
XMCB_2X4<20> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[40] WL[41] S1AHSF400W40_MCB_2X4
XMCB_2X4<21> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[42] WL[43] S1AHSF400W40_MCB_2X4
XMCB_2X4<22> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[44] WL[45] S1AHSF400W40_MCB_2X4
XMCB_2X4<23> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[46] WL[47] S1AHSF400W40_MCB_2X4
XMCB_2X4<24> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[48] WL[49] S1AHSF400W40_MCB_2X4
XMCB_2X4<25> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[50] WL[51] S1AHSF400W40_MCB_2X4
XMCB_2X4<26> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[52] WL[53] S1AHSF400W40_MCB_2X4
XMCB_2X4<27> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[54] WL[55] S1AHSF400W40_MCB_2X4
XMCB_2X4<28> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[56] WL[57] S1AHSF400W40_MCB_2X4
XMCB_2X4<29> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[58] WL[59] S1AHSF400W40_MCB_2X4
XMCB_2X4<30> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[60] WL[61] S1AHSF400W40_MCB_2X4
XMCB_2X4<31> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[62] WL[63] S1AHSF400W40_MCB_2X4
XMCB_2X4<32> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[64] WL[65] S1AHSF400W40_MCB_2X4
XMCB_2X4<33> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[66] WL[67] S1AHSF400W40_MCB_2X4
XMCB_2X4<34> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[68] WL[69] S1AHSF400W40_MCB_2X4
XMCB_2X4<35> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[70] WL[71] S1AHSF400W40_MCB_2X4
XMCB_2X4<36> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[72] WL[73] S1AHSF400W40_MCB_2X4
XMCB_2X4<37> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[74] WL[75] S1AHSF400W40_MCB_2X4
XMCB_2X4<38> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[76] WL[77] S1AHSF400W40_MCB_2X4
XMCB_2X4<39> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[78] WL[79] S1AHSF400W40_MCB_2X4
XMCB_2X4<40> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[80] WL[81] S1AHSF400W40_MCB_2X4
XMCB_2X4<41> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[82] WL[83] S1AHSF400W40_MCB_2X4
XMCB_2X4<42> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[84] WL[85] S1AHSF400W40_MCB_2X4
XMCB_2X4<43> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[86] WL[87] S1AHSF400W40_MCB_2X4
XMCB_2X4<44> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[88] WL[89] S1AHSF400W40_MCB_2X4
XMCB_2X4<45> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[90] WL[91] S1AHSF400W40_MCB_2X4
XMCB_2X4<46> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[92] WL[93] S1AHSF400W40_MCB_2X4
XMCB_2X4<47> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[94] WL[95] S1AHSF400W40_MCB_2X4
XMCB_2X4<48> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[96] WL[97] S1AHSF400W40_MCB_2X4
XMCB_2X4<49> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[98] WL[99] S1AHSF400W40_MCB_2X4
XMCB_2X4<50> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[100] WL[101] S1AHSF400W40_MCB_2X4
XMCB_2X4<51> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[102] WL[103] S1AHSF400W40_MCB_2X4
XMCB_2X4<52> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[104] WL[105] S1AHSF400W40_MCB_2X4
XMCB_2X4<53> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[106] WL[107] S1AHSF400W40_MCB_2X4
XMCB_2X4<54> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[108] WL[109] S1AHSF400W40_MCB_2X4
XMCB_2X4<55> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[110] WL[111] S1AHSF400W40_MCB_2X4
XMCB_2X4<56> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[112] WL[113] S1AHSF400W40_MCB_2X4
XMCB_2X4<57> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[114] WL[115] S1AHSF400W40_MCB_2X4
XMCB_2X4<58> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[116] WL[117] S1AHSF400W40_MCB_2X4
XMCB_2X4<59> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[118] WL[119] S1AHSF400W40_MCB_2X4
XMCB_2X4<60> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[120] WL[121] S1AHSF400W40_MCB_2X4
XMCB_2X4<61> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[122] WL[123] S1AHSF400W40_MCB_2X4
XMCB_2X4<62> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[124] WL[125] S1AHSF400W40_MCB_2X4
XMCB_2X4<63> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[126] WL[127] S1AHSF400W40_MCB_2X4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    MCB_256X4_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_256X4_CHAR BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL 
+ GBLB GW GWB VDDI VSSI WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] 
+ WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] 
+ WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] 
+ WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] 
+ WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] 
+ WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] 
+ WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] WL[72] WL[73] WL[74] 
+ WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] WL[83] WL[84] WL[85] 
+ WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] WL[94] WL[95] WL[96] 
+ WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] WL[104] WL[105] WL[106] 
+ WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] WL[113] WL[114] WL[115] 
+ WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] WL[122] WL[123] WL[124] 
+ WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] WL[131] WL[132] WL[133] 
+ WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] WL[140] WL[141] WL[142] 
+ WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] WL[149] WL[150] WL[151] 
+ WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] WL[158] WL[159] WL[160] 
+ WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] WL[167] WL[168] WL[169] 
+ WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] WL[176] WL[177] WL[178] 
+ WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] WL[185] WL[186] WL[187] 
+ WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] WL[194] WL[195] WL[196] 
+ WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] WL[203] WL[204] WL[205] 
+ WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] WL[212] WL[213] WL[214] 
+ WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] WL[221] WL[222] WL[223] 
+ WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] WL[230] WL[231] WL[232] 
+ WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] WL[239] WL[240] WL[241] 
+ WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] WL[248] WL[249] WL[250] 
+ WL[251] WL[252] WL[253] WL[254] WL[255]
*.PININFO WL[0]:I WL[1]:I WL[2]:I WL[3]:I WL[4]:I WL[5]:I WL[6]:I WL[7]:I 
*.PININFO WL[8]:I WL[9]:I WL[10]:I WL[11]:I WL[12]:I WL[13]:I WL[14]:I 
*.PININFO WL[15]:I WL[16]:I WL[17]:I WL[18]:I WL[19]:I WL[20]:I WL[21]:I 
*.PININFO WL[22]:I WL[23]:I WL[24]:I WL[25]:I WL[26]:I WL[27]:I WL[28]:I 
*.PININFO WL[29]:I WL[30]:I WL[31]:I WL[32]:I WL[33]:I WL[34]:I WL[35]:I 
*.PININFO WL[36]:I WL[37]:I WL[38]:I WL[39]:I WL[40]:I WL[41]:I WL[42]:I 
*.PININFO WL[43]:I WL[44]:I WL[45]:I WL[46]:I WL[47]:I WL[48]:I WL[49]:I 
*.PININFO WL[50]:I WL[51]:I WL[52]:I WL[53]:I WL[54]:I WL[55]:I WL[56]:I 
*.PININFO WL[57]:I WL[58]:I WL[59]:I WL[60]:I WL[61]:I WL[62]:I WL[63]:I 
*.PININFO WL[64]:I WL[65]:I WL[66]:I WL[67]:I WL[68]:I WL[69]:I WL[70]:I 
*.PININFO WL[71]:I WL[72]:I WL[73]:I WL[74]:I WL[75]:I WL[76]:I WL[77]:I 
*.PININFO WL[78]:I WL[79]:I WL[80]:I WL[81]:I WL[82]:I WL[83]:I WL[84]:I 
*.PININFO WL[85]:I WL[86]:I WL[87]:I WL[88]:I WL[89]:I WL[90]:I WL[91]:I 
*.PININFO WL[92]:I WL[93]:I WL[94]:I WL[95]:I WL[96]:I WL[97]:I WL[98]:I 
*.PININFO WL[99]:I WL[100]:I WL[101]:I WL[102]:I WL[103]:I WL[104]:I WL[105]:I 
*.PININFO WL[106]:I WL[107]:I WL[108]:I WL[109]:I WL[110]:I WL[111]:I 
*.PININFO WL[112]:I WL[113]:I WL[114]:I WL[115]:I WL[116]:I WL[117]:I 
*.PININFO WL[118]:I WL[119]:I WL[120]:I WL[121]:I WL[122]:I WL[123]:I 
*.PININFO WL[124]:I WL[125]:I WL[126]:I WL[127]:I WL[128]:I WL[129]:I 
*.PININFO WL[130]:I WL[131]:I WL[132]:I WL[133]:I WL[134]:I WL[135]:I 
*.PININFO WL[136]:I WL[137]:I WL[138]:I WL[139]:I WL[140]:I WL[141]:I 
*.PININFO WL[142]:I WL[143]:I WL[144]:I WL[145]:I WL[146]:I WL[147]:I 
*.PININFO WL[148]:I WL[149]:I WL[150]:I WL[151]:I WL[152]:I WL[153]:I 
*.PININFO WL[154]:I WL[155]:I WL[156]:I WL[157]:I WL[158]:I WL[159]:I 
*.PININFO WL[160]:I WL[161]:I WL[162]:I WL[163]:I WL[164]:I WL[165]:I 
*.PININFO WL[166]:I WL[167]:I WL[168]:I WL[169]:I WL[170]:I WL[171]:I 
*.PININFO WL[172]:I WL[173]:I WL[174]:I WL[175]:I WL[176]:I WL[177]:I 
*.PININFO WL[178]:I WL[179]:I WL[180]:I WL[181]:I WL[182]:I WL[183]:I 
*.PININFO WL[184]:I WL[185]:I WL[186]:I WL[187]:I WL[188]:I WL[189]:I 
*.PININFO WL[190]:I WL[191]:I WL[192]:I WL[193]:I WL[194]:I WL[195]:I 
*.PININFO WL[196]:I WL[197]:I WL[198]:I WL[199]:I WL[200]:I WL[201]:I 
*.PININFO WL[202]:I WL[203]:I WL[204]:I WL[205]:I WL[206]:I WL[207]:I 
*.PININFO WL[208]:I WL[209]:I WL[210]:I WL[211]:I WL[212]:I WL[213]:I 
*.PININFO WL[214]:I WL[215]:I WL[216]:I WL[217]:I WL[218]:I WL[219]:I 
*.PININFO WL[220]:I WL[221]:I WL[222]:I WL[223]:I WL[224]:I WL[225]:I 
*.PININFO WL[226]:I WL[227]:I WL[228]:I WL[229]:I WL[230]:I WL[231]:I 
*.PININFO WL[232]:I WL[233]:I WL[234]:I WL[235]:I WL[236]:I WL[237]:I 
*.PININFO WL[238]:I WL[239]:I WL[240]:I WL[241]:I WL[242]:I WL[243]:I 
*.PININFO WL[244]:I WL[245]:I WL[246]:I WL[247]:I WL[248]:I WL[249]:I 
*.PININFO WL[250]:I WL[251]:I WL[252]:I WL[253]:I WL[254]:I WL[255]:I BL[0]:B 
*.PININFO BL[1]:B BL[2]:B BL[3]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B GBL:B 
*.PININFO GBLB:B GW:B GWB:B VDDI:B VSSI:B
XMCB_2X4<0> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_2X4<1> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[2] WL[3] S1AHSF400W40_MCB_2X4
XMCB_2X4<2> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[4] WL[5] S1AHSF400W40_MCB_2X4
XMCB_2X4<3> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[6] WL[7] S1AHSF400W40_MCB_2X4
XMCB_2X4<4> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[8] WL[9] S1AHSF400W40_MCB_2X4
XMCB_2X4<5> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[10] WL[11] S1AHSF400W40_MCB_2X4
XMCB_2X4<6> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[12] WL[13] S1AHSF400W40_MCB_2X4
XMCB_2X4<7> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[14] WL[15] S1AHSF400W40_MCB_2X4
XMCB_2X4<8> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[16] WL[17] S1AHSF400W40_MCB_2X4
XMCB_2X4<9> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[18] WL[19] S1AHSF400W40_MCB_2X4
XMCB_2X4<10> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[20] WL[21] S1AHSF400W40_MCB_2X4
XMCB_2X4<11> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[22] WL[23] S1AHSF400W40_MCB_2X4
XMCB_2X4<12> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[24] WL[25] S1AHSF400W40_MCB_2X4
XMCB_2X4<13> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[26] WL[27] S1AHSF400W40_MCB_2X4
XMCB_2X4<14> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[28] WL[29] S1AHSF400W40_MCB_2X4
XMCB_2X4<15> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[30] WL[31] S1AHSF400W40_MCB_2X4
XMCB_2X4<16> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[32] WL[33] S1AHSF400W40_MCB_2X4
XMCB_2X4<17> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[34] WL[35] S1AHSF400W40_MCB_2X4
XMCB_2X4<18> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[36] WL[37] S1AHSF400W40_MCB_2X4
XMCB_2X4<19> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[38] WL[39] S1AHSF400W40_MCB_2X4
XMCB_2X4<20> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[40] WL[41] S1AHSF400W40_MCB_2X4
XMCB_2X4<21> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[42] WL[43] S1AHSF400W40_MCB_2X4
XMCB_2X4<22> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[44] WL[45] S1AHSF400W40_MCB_2X4
XMCB_2X4<23> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[46] WL[47] S1AHSF400W40_MCB_2X4
XMCB_2X4<24> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[48] WL[49] S1AHSF400W40_MCB_2X4
XMCB_2X4<25> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[50] WL[51] S1AHSF400W40_MCB_2X4
XMCB_2X4<26> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[52] WL[53] S1AHSF400W40_MCB_2X4
XMCB_2X4<27> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[54] WL[55] S1AHSF400W40_MCB_2X4
XMCB_2X4<28> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[56] WL[57] S1AHSF400W40_MCB_2X4
XMCB_2X4<29> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[58] WL[59] S1AHSF400W40_MCB_2X4
XMCB_2X4<30> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[60] WL[61] S1AHSF400W40_MCB_2X4
XMCB_2X4<31> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[62] WL[63] S1AHSF400W40_MCB_2X4
XMCB_2X4<32> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[64] WL[65] S1AHSF400W40_MCB_2X4
XMCB_2X4<33> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[66] WL[67] S1AHSF400W40_MCB_2X4
XMCB_2X4<34> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[68] WL[69] S1AHSF400W40_MCB_2X4
XMCB_2X4<35> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[70] WL[71] S1AHSF400W40_MCB_2X4
XMCB_2X4<36> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[72] WL[73] S1AHSF400W40_MCB_2X4
XMCB_2X4<37> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[74] WL[75] S1AHSF400W40_MCB_2X4
XMCB_2X4<38> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[76] WL[77] S1AHSF400W40_MCB_2X4
XMCB_2X4<39> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[78] WL[79] S1AHSF400W40_MCB_2X4
XMCB_2X4<40> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[80] WL[81] S1AHSF400W40_MCB_2X4
XMCB_2X4<41> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[82] WL[83] S1AHSF400W40_MCB_2X4
XMCB_2X4<42> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[84] WL[85] S1AHSF400W40_MCB_2X4
XMCB_2X4<43> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[86] WL[87] S1AHSF400W40_MCB_2X4
XMCB_2X4<44> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[88] WL[89] S1AHSF400W40_MCB_2X4
XMCB_2X4<45> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[90] WL[91] S1AHSF400W40_MCB_2X4
XMCB_2X4<46> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[92] WL[93] S1AHSF400W40_MCB_2X4
XMCB_2X4<47> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[94] WL[95] S1AHSF400W40_MCB_2X4
XMCB_2X4<48> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[96] WL[97] S1AHSF400W40_MCB_2X4
XMCB_2X4<49> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[98] WL[99] S1AHSF400W40_MCB_2X4
XMCB_2X4<50> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[100] WL[101] S1AHSF400W40_MCB_2X4
XMCB_2X4<51> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[102] WL[103] S1AHSF400W40_MCB_2X4
XMCB_2X4<52> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[104] WL[105] S1AHSF400W40_MCB_2X4
XMCB_2X4<53> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[106] WL[107] S1AHSF400W40_MCB_2X4
XMCB_2X4<54> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[108] WL[109] S1AHSF400W40_MCB_2X4
XMCB_2X4<55> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[110] WL[111] S1AHSF400W40_MCB_2X4
XMCB_2X4<56> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[112] WL[113] S1AHSF400W40_MCB_2X4
XMCB_2X4<57> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[114] WL[115] S1AHSF400W40_MCB_2X4
XMCB_2X4<58> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[116] WL[117] S1AHSF400W40_MCB_2X4
XMCB_2X4<59> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[118] WL[119] S1AHSF400W40_MCB_2X4
XMCB_2X4<60> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[120] WL[121] S1AHSF400W40_MCB_2X4
XMCB_2X4<61> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[122] WL[123] S1AHSF400W40_MCB_2X4
XMCB_2X4<62> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[124] WL[125] S1AHSF400W40_MCB_2X4
XMCB_2X4<63> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[126] WL[127] S1AHSF400W40_MCB_2X4
XMCB_2X4<64> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[128] WL[129] S1AHSF400W40_MCB_2X4
XMCB_2X4<65> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[130] WL[131] S1AHSF400W40_MCB_2X4
XMCB_2X4<66> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[132] WL[133] S1AHSF400W40_MCB_2X4
XMCB_2X4<67> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[134] WL[135] S1AHSF400W40_MCB_2X4
XMCB_2X4<68> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[136] WL[137] S1AHSF400W40_MCB_2X4
XMCB_2X4<69> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[138] WL[139] S1AHSF400W40_MCB_2X4
XMCB_2X4<70> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[140] WL[141] S1AHSF400W40_MCB_2X4
XMCB_2X4<71> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[142] WL[143] S1AHSF400W40_MCB_2X4
XMCB_2X4<72> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[144] WL[145] S1AHSF400W40_MCB_2X4
XMCB_2X4<73> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[146] WL[147] S1AHSF400W40_MCB_2X4
XMCB_2X4<74> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[148] WL[149] S1AHSF400W40_MCB_2X4
XMCB_2X4<75> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[150] WL[151] S1AHSF400W40_MCB_2X4
XMCB_2X4<76> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[152] WL[153] S1AHSF400W40_MCB_2X4
XMCB_2X4<77> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[154] WL[155] S1AHSF400W40_MCB_2X4
XMCB_2X4<78> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[156] WL[157] S1AHSF400W40_MCB_2X4
XMCB_2X4<79> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[158] WL[159] S1AHSF400W40_MCB_2X4
XMCB_2X4<80> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[160] WL[161] S1AHSF400W40_MCB_2X4
XMCB_2X4<81> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[162] WL[163] S1AHSF400W40_MCB_2X4
XMCB_2X4<82> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[164] WL[165] S1AHSF400W40_MCB_2X4
XMCB_2X4<83> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[166] WL[167] S1AHSF400W40_MCB_2X4
XMCB_2X4<84> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[168] WL[169] S1AHSF400W40_MCB_2X4
XMCB_2X4<85> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[170] WL[171] S1AHSF400W40_MCB_2X4
XMCB_2X4<86> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[172] WL[173] S1AHSF400W40_MCB_2X4
XMCB_2X4<87> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[174] WL[175] S1AHSF400W40_MCB_2X4
XMCB_2X4<88> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[176] WL[177] S1AHSF400W40_MCB_2X4
XMCB_2X4<89> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[178] WL[179] S1AHSF400W40_MCB_2X4
XMCB_2X4<90> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[180] WL[181] S1AHSF400W40_MCB_2X4
XMCB_2X4<91> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[182] WL[183] S1AHSF400W40_MCB_2X4
XMCB_2X4<92> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[184] WL[185] S1AHSF400W40_MCB_2X4
XMCB_2X4<93> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[186] WL[187] S1AHSF400W40_MCB_2X4
XMCB_2X4<94> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[188] WL[189] S1AHSF400W40_MCB_2X4
XMCB_2X4<95> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[190] WL[191] S1AHSF400W40_MCB_2X4
XMCB_2X4<96> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[192] WL[193] S1AHSF400W40_MCB_2X4
XMCB_2X4<97> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[194] WL[195] S1AHSF400W40_MCB_2X4
XMCB_2X4<98> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[196] WL[197] S1AHSF400W40_MCB_2X4
XMCB_2X4<99> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[198] WL[199] S1AHSF400W40_MCB_2X4
XMCB_2X4<100> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[200] WL[201] S1AHSF400W40_MCB_2X4
XMCB_2X4<101> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[202] WL[203] S1AHSF400W40_MCB_2X4
XMCB_2X4<102> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[204] WL[205] S1AHSF400W40_MCB_2X4
XMCB_2X4<103> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[206] WL[207] S1AHSF400W40_MCB_2X4
XMCB_2X4<104> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[208] WL[209] S1AHSF400W40_MCB_2X4
XMCB_2X4<105> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[210] WL[211] S1AHSF400W40_MCB_2X4
XMCB_2X4<106> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[212] WL[213] S1AHSF400W40_MCB_2X4
XMCB_2X4<107> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[214] WL[215] S1AHSF400W40_MCB_2X4
XMCB_2X4<108> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[216] WL[217] S1AHSF400W40_MCB_2X4
XMCB_2X4<109> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[218] WL[219] S1AHSF400W40_MCB_2X4
XMCB_2X4<110> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[220] WL[221] S1AHSF400W40_MCB_2X4
XMCB_2X4<111> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[222] WL[223] S1AHSF400W40_MCB_2X4
XMCB_2X4<112> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[224] WL[225] S1AHSF400W40_MCB_2X4
XMCB_2X4<113> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[226] WL[227] S1AHSF400W40_MCB_2X4
XMCB_2X4<114> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[228] WL[229] S1AHSF400W40_MCB_2X4
XMCB_2X4<115> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[230] WL[231] S1AHSF400W40_MCB_2X4
XMCB_2X4<116> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[232] WL[233] S1AHSF400W40_MCB_2X4
XMCB_2X4<117> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[234] WL[235] S1AHSF400W40_MCB_2X4
XMCB_2X4<118> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[236] WL[237] S1AHSF400W40_MCB_2X4
XMCB_2X4<119> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[238] WL[239] S1AHSF400W40_MCB_2X4
XMCB_2X4<120> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[240] WL[241] S1AHSF400W40_MCB_2X4
XMCB_2X4<121> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[242] WL[243] S1AHSF400W40_MCB_2X4
XMCB_2X4<122> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[244] WL[245] S1AHSF400W40_MCB_2X4
XMCB_2X4<123> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[246] WL[247] S1AHSF400W40_MCB_2X4
XMCB_2X4<124> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[248] WL[249] S1AHSF400W40_MCB_2X4
XMCB_2X4<125> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[250] WL[251] S1AHSF400W40_MCB_2X4
XMCB_2X4<126> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[252] WL[253] S1AHSF400W40_MCB_2X4
XMCB_2X4<127> BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL GBLB GW 
+ GWB VDDI VSSI WL[254] WL[255] S1AHSF400W40_MCB_2X4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    ARR_BLLD_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ARR_BLLD_SIM BLB_BT[0] BLB_BT[1] BLB_TP[0] BLB_TP[1] BL_BT[0] BL_BT[1] 
+ BL_TP[0] BL_TP[1] CVDDI GBLB_BT GBLB_TP GBL_BT GBL_TP GWB_BT GWB_TP GW_BT 
+ GW_TP VDDHD VDDI VSSI
*.PININFO BLB_BT[0]:B BLB_BT[1]:B BLB_TP[0]:B BLB_TP[1]:B BL_BT[0]:B 
*.PININFO BL_BT[1]:B BL_TP[0]:B BL_TP[1]:B CVDDI:B GBLB_BT:B GBLB_TP:B 
*.PININFO GBL_BT:B GBL_TP:B GWB_BT:B GWB_TP:B GW_BT:B GW_TP:B VDDHD:B VDDI:B 
*.PININFO VSSI:B
XI33 NET23[0] NET23[1] NET23[2] NET23[3] NET17[0] NET17[1] NET17[2] NET17[3] 
+ NET24 NET19 NET20 NET18 NET22 NET21 NET017[0] NET017[1] NET017[2] NET017[3] 
+ NET017[4] NET017[5] NET017[6] NET017[7] NET017[8] NET017[9] NET017[10] 
+ NET017[11] NET017[12] NET017[13] NET017[14] NET017[15] NET017[16] NET017[17] 
+ NET017[18] NET017[19] NET017[20] NET017[21] NET017[22] NET017[23] NET017[24] 
+ NET017[25] NET017[26] NET017[27] NET017[28] NET017[29] NET017[30] NET017[31] 
+ S1AHSF400W40_MCB_32X4_CHAR
XI34 NET030[0] NET030[1] NET030[2] NET030[3] NET029[0] NET029[1] NET029[2] 
+ NET029[3] NET034 NET033 NET027 NET028 NET031 NET032 NET026[0] NET026[1] 
+ NET026[2] NET026[3] NET026[4] NET026[5] NET026[6] NET026[7] NET026[8] 
+ NET026[9] NET026[10] NET026[11] NET026[12] NET026[13] NET026[14] NET026[15] 
+ NET026[16] NET026[17] NET026[18] NET026[19] NET026[20] NET026[21] NET026[22] 
+ NET026[23] NET026[24] NET026[25] NET026[26] NET026[27] NET026[28] NET026[29] 
+ NET026[30] NET026[31] NET026[32] NET026[33] NET026[34] NET026[35] NET026[36] 
+ NET026[37] NET026[38] NET026[39] NET026[40] NET026[41] NET026[42] NET026[43] 
+ NET026[44] NET026[45] NET026[46] NET026[47] NET026[48] NET026[49] NET026[50] 
+ NET026[51] NET026[52] NET026[53] NET026[54] NET026[55] NET026[56] NET026[57] 
+ NET026[58] NET026[59] NET026[60] NET026[61] NET026[62] NET026[63] 
+ S1AHSF400W40_MCB_64X4_CHAR
XI35 NET039[0] NET039[1] NET039[2] NET039[3] NET038[0] NET038[1] NET038[2] 
+ NET038[3] NET043 NET042 NET036 NET037 NET040 NET041 NET035[0] NET035[1] 
+ NET035[2] NET035[3] NET035[4] NET035[5] NET035[6] NET035[7] NET035[8] 
+ NET035[9] NET035[10] NET035[11] NET035[12] NET035[13] NET035[14] NET035[15] 
+ NET035[16] NET035[17] NET035[18] NET035[19] NET035[20] NET035[21] NET035[22] 
+ NET035[23] NET035[24] NET035[25] NET035[26] NET035[27] NET035[28] NET035[29] 
+ NET035[30] NET035[31] NET035[32] NET035[33] NET035[34] NET035[35] NET035[36] 
+ NET035[37] NET035[38] NET035[39] NET035[40] NET035[41] NET035[42] NET035[43] 
+ NET035[44] NET035[45] NET035[46] NET035[47] NET035[48] NET035[49] NET035[50] 
+ NET035[51] NET035[52] NET035[53] NET035[54] NET035[55] NET035[56] NET035[57] 
+ NET035[58] NET035[59] NET035[60] NET035[61] NET035[62] NET035[63] NET035[64] 
+ NET035[65] NET035[66] NET035[67] NET035[68] NET035[69] NET035[70] NET035[71] 
+ NET035[72] NET035[73] NET035[74] NET035[75] NET035[76] NET035[77] NET035[78] 
+ NET035[79] NET035[80] NET035[81] NET035[82] NET035[83] NET035[84] NET035[85] 
+ NET035[86] NET035[87] NET035[88] NET035[89] NET035[90] NET035[91] NET035[92] 
+ NET035[93] NET035[94] NET035[95] NET035[96] NET035[97] NET035[98] NET035[99] 
+ NET035[100] NET035[101] NET035[102] NET035[103] NET035[104] NET035[105] 
+ NET035[106] NET035[107] NET035[108] NET035[109] NET035[110] NET035[111] 
+ NET035[112] NET035[113] NET035[114] NET035[115] NET035[116] NET035[117] 
+ NET035[118] NET035[119] NET035[120] NET035[121] NET035[122] NET035[123] 
+ NET035[124] NET035[125] NET035[126] NET035[127] S1AHSF400W40_MCB_128X4_CHAR
XI36 NET048[0] NET048[1] NET048[2] NET048[3] NET047[0] NET047[1] NET047[2] 
+ NET047[3] NET052 NET051 NET045 NET046 NET049 NET050 NET044[0] NET044[1] 
+ NET044[2] NET044[3] NET044[4] NET044[5] NET044[6] NET044[7] NET044[8] 
+ NET044[9] NET044[10] NET044[11] NET044[12] NET044[13] NET044[14] NET044[15] 
+ NET044[16] NET044[17] NET044[18] NET044[19] NET044[20] NET044[21] NET044[22] 
+ NET044[23] NET044[24] NET044[25] NET044[26] NET044[27] NET044[28] NET044[29] 
+ NET044[30] NET044[31] NET044[32] NET044[33] NET044[34] NET044[35] NET044[36] 
+ NET044[37] NET044[38] NET044[39] NET044[40] NET044[41] NET044[42] NET044[43] 
+ NET044[44] NET044[45] NET044[46] NET044[47] NET044[48] NET044[49] NET044[50] 
+ NET044[51] NET044[52] NET044[53] NET044[54] NET044[55] NET044[56] NET044[57] 
+ NET044[58] NET044[59] NET044[60] NET044[61] NET044[62] NET044[63] NET044[64] 
+ NET044[65] NET044[66] NET044[67] NET044[68] NET044[69] NET044[70] NET044[71] 
+ NET044[72] NET044[73] NET044[74] NET044[75] NET044[76] NET044[77] NET044[78] 
+ NET044[79] NET044[80] NET044[81] NET044[82] NET044[83] NET044[84] NET044[85] 
+ NET044[86] NET044[87] NET044[88] NET044[89] NET044[90] NET044[91] NET044[92] 
+ NET044[93] NET044[94] NET044[95] NET044[96] NET044[97] NET044[98] NET044[99] 
+ NET044[100] NET044[101] NET044[102] NET044[103] NET044[104] NET044[105] 
+ NET044[106] NET044[107] NET044[108] NET044[109] NET044[110] NET044[111] 
+ NET044[112] NET044[113] NET044[114] NET044[115] NET044[116] NET044[117] 
+ NET044[118] NET044[119] NET044[120] NET044[121] NET044[122] NET044[123] 
+ NET044[124] NET044[125] NET044[126] NET044[127] NET044[128] NET044[129] 
+ NET044[130] NET044[131] NET044[132] NET044[133] NET044[134] NET044[135] 
+ NET044[136] NET044[137] NET044[138] NET044[139] NET044[140] NET044[141] 
+ NET044[142] NET044[143] NET044[144] NET044[145] NET044[146] NET044[147] 
+ NET044[148] NET044[149] NET044[150] NET044[151] NET044[152] NET044[153] 
+ NET044[154] NET044[155] NET044[156] NET044[157] NET044[158] NET044[159] 
+ NET044[160] NET044[161] NET044[162] NET044[163] NET044[164] NET044[165] 
+ NET044[166] NET044[167] NET044[168] NET044[169] NET044[170] NET044[171] 
+ NET044[172] NET044[173] NET044[174] NET044[175] NET044[176] NET044[177] 
+ NET044[178] NET044[179] NET044[180] NET044[181] NET044[182] NET044[183] 
+ NET044[184] NET044[185] NET044[186] NET044[187] NET044[188] NET044[189] 
+ NET044[190] NET044[191] NET044[192] NET044[193] NET044[194] NET044[195] 
+ NET044[196] NET044[197] NET044[198] NET044[199] NET044[200] NET044[201] 
+ NET044[202] NET044[203] NET044[204] NET044[205] NET044[206] NET044[207] 
+ NET044[208] NET044[209] NET044[210] NET044[211] NET044[212] NET044[213] 
+ NET044[214] NET044[215] NET044[216] NET044[217] NET044[218] NET044[219] 
+ NET044[220] NET044[221] NET044[222] NET044[223] NET044[224] NET044[225] 
+ NET044[226] NET044[227] NET044[228] NET044[229] NET044[230] NET044[231] 
+ NET044[232] NET044[233] NET044[234] NET044[235] NET044[236] NET044[237] 
+ NET044[238] NET044[239] NET044[240] NET044[241] NET044[242] NET044[243] 
+ NET044[244] NET044[245] NET044[246] NET044[247] NET044[248] NET044[249] 
+ NET044[250] NET044[251] NET044[252] NET044[253] NET044[254] NET044[255] 
+ S1AHSF400W40_MCB_256X4_CHAR
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    MCB_2X4_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_2X4_CHAR BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL 
+ GBLB GW GWB VDDI VSSI WL[0] WL[1]
*.PININFO WL[0]:I WL[1]:I BL[0]:B BL[1]:B BL[2]:B BL[3]:B BLB[0]:B BLB[1]:B 
*.PININFO BLB[2]:B BLB[3]:B GBL:B GBLB:B GW:B GWB:B VDDI:B VSSI:B
XMCB_0<0> BL[0] BLB[0] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<1> BL[1] BLB[1] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<2> BL[2] BLB[2] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<3> BL[3] BLB[3] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_1<0> BL[0] BLB[0] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<1> BL[1] BLB[1] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<2> BL[2] BLB[2] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<3> BL[3] BLB[3] VDDI VSSI WL[1] S1AHSF400W40_MCB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    ARR_WLLD_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ARR_WLLD_SIM CVDDI VDDHD VDDI VSSI WL_LT[0] WL_LT[1] WL_RT[0] WL_RT[1]
*.PININFO CVDDI:B VDDHD:B VDDI:B VSSI:B WL_LT[0]:B WL_LT[1]:B WL_RT[0]:B 
*.PININFO WL_RT[1]:B
XI21 NET011[0] NET011[1] NET011[2] NET011[3] NET07[0] NET07[1] NET07[2] 
+ NET07[3] NET014 NET012 NET013 NET01 NET11 NET10 NET04[0] NET04[1] 
+ S1AHSF400W40_MCB_2X4_CHAR
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    ARR_MCB_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ARR_MCB_SIM BL[0] BL[1] BLB[0] BLB[1] CVDDI GBL GBLB GW GWB VDDHD VDDI 
+ VSSI WL_LT[0] WL_LT[1] WL_RT[0] WL_RT[1]
*.PININFO BL[0]:B BL[1]:B BLB[0]:B BLB[1]:B CVDDI:B GBL:B GBLB:B GW:B GWB:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WL_LT[0]:B WL_LT[1]:B WL_RT[0]:B WL_RT[1]:B
XI22 NET021[0] NET021[1] NET021[2] NET021[3] NET01[0] NET01[1] NET01[2] 
+ NET01[3] NET022 NET017 NET018 NET02 NET020 NET019 NET03[0] NET03[1] 
+ S1AHSF400W40_MCB_2X4_CHAR
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    PRECHARGE
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_PRECHARGE BL BLB BLEQB VDDI
*.PININFO BLEQB:I BL:B BLB:B VDDI:B
MP17 BLB BLEQB VDDI VDDI PCH L=60N W=800N M=2
MP5 BL BLEQB BLB VDDI PCH L=60N W=800N M=1
MP0 VDDI BLEQB BL VDDI PCH L=60N W=800N M=2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    YPASS_M8
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_YPASS_M8 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BLB[0] BLB[1] 
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLEQ BLEQB DL DLB READ VDDI VSSI 
+ WC WRITE WT Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7]
*.PININFO BLEQ:I READ:I WRITE:I Y[0]:I Y[1]:I Y[2]:I Y[3]:I Y[4]:I Y[5]:I 
*.PININFO Y[6]:I Y[7]:I BLEQB:O BL[0]:B BL[1]:B BL[2]:B BL[3]:B BL[4]:B 
*.PININFO BL[5]:B BL[6]:B BL[7]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B BLB[4]:B 
*.PININFO BLB[5]:B BLB[6]:B BLB[7]:B DL:B DLB:B VDDI:B VSSI:B WC:B WT:B
XPRECHARGE<0> BL[0] BLB[0] BLEQB VDDI S1AHSF400W40_PRECHARGE
XPRECHARGE<1> BL[1] BLB[1] BLEQB VDDI S1AHSF400W40_PRECHARGE
XPRECHARGE<2> BL[2] BLB[2] BLEQB VDDI S1AHSF400W40_PRECHARGE
XPRECHARGE<3> BL[3] BLB[3] BLEQB VDDI S1AHSF400W40_PRECHARGE
XPRECHARGE<4> BL[4] BLB[4] BLEQB VDDI S1AHSF400W40_PRECHARGE
XPRECHARGE<5> BL[5] BLB[5] BLEQB VDDI S1AHSF400W40_PRECHARGE
XPRECHARGE<6> BL[6] BLB[6] BLEQB VDDI S1AHSF400W40_PRECHARGE
XPRECHARGE<7> BL[7] BLB[7] BLEQB VDDI S1AHSF400W40_PRECHARGE
XI252<0> Y[0] NET0112[0] VSSI VDDI VDDI YB_WRITE[0] S1AHSF400W40_INV_BULK FN=1 WN=0.36U 
+ LN=0.06U FP=1 WP=0.36U LP=0.06U M=1
XI252<1> Y[1] NET0112[1] VSSI VDDI VDDI YB_WRITE[1] S1AHSF400W40_INV_BULK FN=1 WN=0.36U 
+ LN=0.06U FP=1 WP=0.36U LP=0.06U M=1
XI252<2> Y[2] NET0112[2] VSSI VDDI VDDI YB_WRITE[2] S1AHSF400W40_INV_BULK FN=1 WN=0.36U 
+ LN=0.06U FP=1 WP=0.36U LP=0.06U M=1
XI252<3> Y[3] NET0112[3] VSSI VDDI VDDI YB_WRITE[3] S1AHSF400W40_INV_BULK FN=1 WN=0.36U 
+ LN=0.06U FP=1 WP=0.36U LP=0.06U M=1
XI252<4> Y[4] NET0112[4] VSSI VDDI VDDI YB_WRITE[4] S1AHSF400W40_INV_BULK FN=1 WN=0.36U 
+ LN=0.06U FP=1 WP=0.36U LP=0.06U M=1
XI252<5> Y[5] NET0112[5] VSSI VDDI VDDI YB_WRITE[5] S1AHSF400W40_INV_BULK FN=1 WN=0.36U 
+ LN=0.06U FP=1 WP=0.36U LP=0.06U M=1
XI252<6> Y[6] NET0112[6] VSSI VDDI VDDI YB_WRITE[6] S1AHSF400W40_INV_BULK FN=1 WN=0.36U 
+ LN=0.06U FP=1 WP=0.36U LP=0.06U M=1
XI252<7> Y[7] NET0112[7] VSSI VDDI VDDI YB_WRITE[7] S1AHSF400W40_INV_BULK FN=1 WN=0.36U 
+ LN=0.06U FP=1 WP=0.36U LP=0.06U M=1
XI249<0> Y[0] NET0116[0] VSSI VDDI VDDI YB_READ[0] S1AHSF400W40_INV_BULK FN=1 WN=0.36U 
+ LN=0.06U FP=1 WP=0.36U LP=0.06U M=1
XI249<1> Y[1] NET0116[1] VSSI VDDI VDDI YB_READ[1] S1AHSF400W40_INV_BULK FN=1 WN=0.36U 
+ LN=0.06U FP=1 WP=0.36U LP=0.06U M=1
XI249<2> Y[2] NET0116[2] VSSI VDDI VDDI YB_READ[2] S1AHSF400W40_INV_BULK FN=1 WN=0.36U 
+ LN=0.06U FP=1 WP=0.36U LP=0.06U M=1
XI249<3> Y[3] NET0116[3] VSSI VDDI VDDI YB_READ[3] S1AHSF400W40_INV_BULK FN=1 WN=0.36U 
+ LN=0.06U FP=1 WP=0.36U LP=0.06U M=1
XI249<4> Y[4] NET0116[4] VSSI VDDI VDDI YB_READ[4] S1AHSF400W40_INV_BULK FN=1 WN=0.36U 
+ LN=0.06U FP=1 WP=0.36U LP=0.06U M=1
XI249<5> Y[5] NET0116[5] VSSI VDDI VDDI YB_READ[5] S1AHSF400W40_INV_BULK FN=1 WN=0.36U 
+ LN=0.06U FP=1 WP=0.36U LP=0.06U M=1
XI249<6> Y[6] NET0116[6] VSSI VDDI VDDI YB_READ[6] S1AHSF400W40_INV_BULK FN=1 WN=0.36U 
+ LN=0.06U FP=1 WP=0.36U LP=0.06U M=1
XI249<7> Y[7] NET0116[7] VSSI VDDI VDDI YB_READ[7] S1AHSF400W40_INV_BULK FN=1 WN=0.36U 
+ LN=0.06U FP=1 WP=0.36U LP=0.06U M=1
MP29<0> YB_WRITE[0] WRITE VDDI VDDI PCH L=60N W=360.0N M=1
MP29<1> YB_WRITE[1] WRITE VDDI VDDI PCH L=60N W=360.0N M=1
MP29<2> YB_WRITE[2] WRITE VDDI VDDI PCH L=60N W=360.0N M=1
MP29<3> YB_WRITE[3] WRITE VDDI VDDI PCH L=60N W=360.0N M=1
MP29<4> YB_WRITE[4] WRITE VDDI VDDI PCH L=60N W=360.0N M=1
MP29<5> YB_WRITE[5] WRITE VDDI VDDI PCH L=60N W=360.0N M=1
MP29<6> YB_WRITE[6] WRITE VDDI VDDI PCH L=60N W=360.0N M=1
MP29<7> YB_WRITE[7] WRITE VDDI VDDI PCH L=60N W=360.0N M=1
MP22 VDDI BLEQB DL VDDI PCH L=60N W=200N M=1
MP0<0> DL YB_READ[0] BL[0] VDDI PCH L=60N W=800N M=1
MP0<1> DL YB_READ[1] BL[1] VDDI PCH L=60N W=800N M=1
MP0<2> DL YB_READ[2] BL[2] VDDI PCH L=60N W=800N M=1
MP0<3> DL YB_READ[3] BL[3] VDDI PCH L=60N W=800N M=1
MP0<4> DL YB_READ[4] BL[4] VDDI PCH L=60N W=800N M=1
MP0<5> DL YB_READ[5] BL[5] VDDI PCH L=60N W=800N M=1
MP0<6> DL YB_READ[6] BL[6] VDDI PCH L=60N W=800N M=1
MP0<7> DL YB_READ[7] BL[7] VDDI PCH L=60N W=800N M=1
MP3 DLB BLEQB VDDI VDDI PCH L=60N W=200N M=1
MP10<0> DLB YB_READ[0] BLB[0] VDDI PCH L=60N W=800N M=1
MP10<1> DLB YB_READ[1] BLB[1] VDDI PCH L=60N W=800N M=1
MP10<2> DLB YB_READ[2] BLB[2] VDDI PCH L=60N W=800N M=1
MP10<3> DLB YB_READ[3] BLB[3] VDDI PCH L=60N W=800N M=1
MP10<4> DLB YB_READ[4] BLB[4] VDDI PCH L=60N W=800N M=1
MP10<5> DLB YB_READ[5] BLB[5] VDDI PCH L=60N W=800N M=1
MP10<6> DLB YB_READ[6] BLB[6] VDDI PCH L=60N W=800N M=1
MP10<7> DLB YB_READ[7] BLB[7] VDDI PCH L=60N W=800N M=1
MP17<0> YB_READ[0] READ VDDI VDDI PCH L=60N W=360.0N M=1
MP17<1> YB_READ[1] READ VDDI VDDI PCH L=60N W=360.0N M=1
MP17<2> YB_READ[2] READ VDDI VDDI PCH L=60N W=360.0N M=1
MP17<3> YB_READ[3] READ VDDI VDDI PCH L=60N W=360.0N M=1
MP17<4> YB_READ[4] READ VDDI VDDI PCH L=60N W=360.0N M=1
MP17<5> YB_READ[5] READ VDDI VDDI PCH L=60N W=360.0N M=1
MP17<6> YB_READ[6] READ VDDI VDDI PCH L=60N W=360.0N M=1
MP17<7> YB_READ[7] READ VDDI VDDI PCH L=60N W=360.0N M=1
MN1<0> NET0112[0] WRITE VSSI VSSI NCH L=60N W=360.0N M=1
MN1<1> NET0112[1] WRITE VSSI VSSI NCH L=60N W=360.0N M=1
MN1<2> NET0112[2] WRITE VSSI VSSI NCH L=60N W=360.0N M=1
MN1<3> NET0112[3] WRITE VSSI VSSI NCH L=60N W=360.0N M=1
MN1<4> NET0112[4] WRITE VSSI VSSI NCH L=60N W=360.0N M=1
MN1<5> NET0112[5] WRITE VSSI VSSI NCH L=60N W=360.0N M=1
MN1<6> NET0112[6] WRITE VSSI VSSI NCH L=60N W=360.0N M=1
MN1<7> NET0112[7] WRITE VSSI VSSI NCH L=60N W=360.0N M=1
MN13<0> NET0116[0] READ VSSI VSSI NCH L=60N W=360.0N M=1
MN13<1> NET0116[1] READ VSSI VSSI NCH L=60N W=360.0N M=1
MN13<2> NET0116[2] READ VSSI VSSI NCH L=60N W=360.0N M=1
MN13<3> NET0116[3] READ VSSI VSSI NCH L=60N W=360.0N M=1
MN13<4> NET0116[4] READ VSSI VSSI NCH L=60N W=360.0N M=1
MN13<5> NET0116[5] READ VSSI VSSI NCH L=60N W=360.0N M=1
MN13<6> NET0116[6] READ VSSI VSSI NCH L=60N W=360.0N M=1
MN13<7> NET0116[7] READ VSSI VSSI NCH L=60N W=360.0N M=1
MN18<0> BLB[0] Y_WRITE[0] WC VSSI NCH L=60N W=1.6U M=1
MN18<1> BLB[1] Y_WRITE[1] WC VSSI NCH L=60N W=1.6U M=1
MN18<2> BLB[2] Y_WRITE[2] WC VSSI NCH L=60N W=1.6U M=1
MN18<3> BLB[3] Y_WRITE[3] WC VSSI NCH L=60N W=1.6U M=1
MN18<4> BLB[4] Y_WRITE[4] WC VSSI NCH L=60N W=1.6U M=1
MN18<5> BLB[5] Y_WRITE[5] WC VSSI NCH L=60N W=1.6U M=1
MN18<6> BLB[6] Y_WRITE[6] WC VSSI NCH L=60N W=1.6U M=1
MN18<7> BLB[7] Y_WRITE[7] WC VSSI NCH L=60N W=1.6U M=1
MN31<0> BL[0] Y_WRITE[0] WT VSSI NCH L=60N W=1.6U M=1
MN31<1> BL[1] Y_WRITE[1] WT VSSI NCH L=60N W=1.6U M=1
MN31<2> BL[2] Y_WRITE[2] WT VSSI NCH L=60N W=1.6U M=1
MN31<3> BL[3] Y_WRITE[3] WT VSSI NCH L=60N W=1.6U M=1
MN31<4> BL[4] Y_WRITE[4] WT VSSI NCH L=60N W=1.6U M=1
MN31<5> BL[5] Y_WRITE[5] WT VSSI NCH L=60N W=1.6U M=1
MN31<6> BL[6] Y_WRITE[6] WT VSSI NCH L=60N W=1.6U M=1
MN31<7> BL[7] Y_WRITE[7] WT VSSI NCH L=60N W=1.6U M=1
XINV0 BLEQ VSSI VDDI BLEQB S1AHSF400W40_AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=1.6U LP=0.06U 
+ M=2
XI214<0> YB_WRITE[0] VSSI VDDI Y_WRITE[0] S1AHSF400W40_AINV FN=1 WN=0.18U LN=0.06U FP=1 
+ WP=0.36U LP=0.06U M=1
XI214<1> YB_WRITE[1] VSSI VDDI Y_WRITE[1] S1AHSF400W40_AINV FN=1 WN=0.18U LN=0.06U FP=1 
+ WP=0.36U LP=0.06U M=1
XI214<2> YB_WRITE[2] VSSI VDDI Y_WRITE[2] S1AHSF400W40_AINV FN=1 WN=0.18U LN=0.06U FP=1 
+ WP=0.36U LP=0.06U M=1
XI214<3> YB_WRITE[3] VSSI VDDI Y_WRITE[3] S1AHSF400W40_AINV FN=1 WN=0.18U LN=0.06U FP=1 
+ WP=0.36U LP=0.06U M=1
XI214<4> YB_WRITE[4] VSSI VDDI Y_WRITE[4] S1AHSF400W40_AINV FN=1 WN=0.18U LN=0.06U FP=1 
+ WP=0.36U LP=0.06U M=1
XI214<5> YB_WRITE[5] VSSI VDDI Y_WRITE[5] S1AHSF400W40_AINV FN=1 WN=0.18U LN=0.06U FP=1 
+ WP=0.36U LP=0.06U M=1
XI214<6> YB_WRITE[6] VSSI VDDI Y_WRITE[6] S1AHSF400W40_AINV FN=1 WN=0.18U LN=0.06U FP=1 
+ WP=0.36U LP=0.06U M=1
XI214<7> YB_WRITE[7] VSSI VDDI Y_WRITE[7] S1AHSF400W40_AINV FN=1 WN=0.18U LN=0.06U FP=1 
+ WP=0.36U LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    SA_M16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SA_M16 DLB_DN_0 DLB_DN_1 DLB_UP_0 DLB_UP_1 DL_DN_0 DL_DN_1 DL_UP_0 
+ DL_UP_1 GBL GBLB PGB_DN_0 PGB_DN_1 PGB_UP_0 PGB_UP_1 PREB SAE VDDI VSSI
*.PININFO PGB_DN_0:I PGB_DN_1:I PGB_UP_0:I PGB_UP_1:I PREB:I SAE:I DLB_DN_0:B 
*.PININFO DLB_DN_1:B DLB_UP_0:B DLB_UP_1:B DL_DN_0:B DL_DN_1:B DL_UP_0:B 
*.PININFO DL_UP_1:B GBL:B GBLB:B VDDI:B VSSI:B
MM6 DL_UP_1 PGB_UP_1 DL_IN VDDI PCH L=100N W=1U M=1
MM5 DLB_IN PGB_UP_0 DLB_UP_0 VDDI PCH L=100N W=1U M=1
MP11 DLB_IN PREB VDDI VDDI PCH L=100N W=1U M=1
MM4 DLB_IN PGB_UP_1 DLB_UP_1 VDDI PCH L=100N W=1U M=1
MM7 DL_UP_0 PGB_UP_0 DL_IN VDDI PCH L=100N W=1U M=1
MP8 DL_IN PREB DLB_IN VDDI PCH L=120.0N W=1U M=2
MP3 DLB_IN DL_IN VDDI VDDI PCH L=120.0N W=1U M=1
MP7 DLB_IN PGB_DN_1 DLB_DN_1 VDDI PCH L=100N W=1U M=1
MP2 VDDI DLB_IN DL_IN VDDI PCH L=120.0N W=1U M=1
MP13 DL_DN_0 PGB_DN_0 DL_IN VDDI PCH L=100N W=1U M=1
MP6 DL_DN_1 PGB_DN_1 DL_IN VDDI PCH L=100N W=1U M=1
MP14 DLB_IN PGB_DN_0 DLB_DN_0 VDDI PCH L=100N W=1U M=1
MP10 DL_IN PREB VDDI VDDI PCH L=100N W=1U M=1
MN12 GBLB SOB VSSI VSSI NCH L=65.0N W=800N M=6
MN11 GBL SO VSSI VSSI NCH L=65.0N W=800N M=6
MN1 DLB_IN DL_IN NS VSSI NCH L=180.0N W=500N M=4
MN2 NS SAE VSSI VSSI NCH L=80N W=500N M=4
MN0 NS DLB_IN DL_IN VSSI NCH L=180.0N W=500N M=4
XINV0 DL_IN VSSI VDDI SO S1AHSF400W40_AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=1U LP=0.06U M=1
XINV1 DLB_IN VSSI VDDI SOB S1AHSF400W40_AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=1U LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    IO_RWBLK_M16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_IO_RWBLK_M16 BLEQB_DN_0 BLEQB_DN_1 BLEQB_UP_0 BLEQB_UP_1 BLEQ_DN 
+ BLEQ_UP DLB_DN_0 DLB_DN_1 DLB_UP_0 DLB_UP_1 DL_DN_0 DL_DN_1 DL_UP_0 DL_UP_1 
+ GBL GBLB GW GWB RE READ SAEB VDDHD VDDI VSSI WC[0] WC[1] WE WRITE WT[0] 
+ WT[1] YL[0] YL[1]
*.PININFO BLEQB_DN_0:I BLEQB_DN_1:I BLEQB_UP_0:I BLEQB_UP_1:I BLEQ_DN:I 
*.PININFO BLEQ_UP:I GW:I GWB:I RE:I SAEB:I WE:I YL[0]:I YL[1]:I READ:O WC[0]:O 
*.PININFO WC[1]:O WRITE:O WT[0]:O WT[1]:O DLB_DN_0:B DLB_DN_1:B DLB_UP_0:B 
*.PININFO DLB_UP_1:B DL_DN_0:B DL_DN_1:B DL_UP_0:B DL_UP_1:B GBL:B GBLB:B 
*.PININFO VDDHD:B VDDI:B VSSI:B
XSA DLB_DN_0 DLB_DN_1 DLB_UP_0 DLB_UP_1 DL_DN_0 DL_DN_1 DL_UP_0 DL_UP_1 GBL 
+ GBLB PGB_DN_0 PGB_DN_1 PGB_UP_0 PGB_UP_1 PREB SAE VDDI VSSI S1AHSF400W40_SA_M16
XI222 SAEC BLEQ_UP BLEQ_DN VSSI VDDI PREB S1AHSF400W40_ANAND3 FN3=1 WN3=0.4U LN3=0.06U 
+ FN2=1 WN2=0.4U LN2=0.06U FN1=1 WN1=0.4U LN1=0.06U FP1=1 WP1=0.4U LP1=0.06U 
+ FP2=1 WP2=0.4U LP2=0.06U FP3=1 WP3=0.4U LP3=0.06U M=1
MM26 LWDC[1] GWDC_YL VDDHD VDDI PCH L=60N W=1U M=1
MM25 GWDC_YL GWB VDDHD VDDI PCH L=60N W=300N M=1
MM31 GWDC_YLB GWB VDDHD VDDI PCH L=60N W=300N M=1
MM30 LWDC[0] GWDC_YLB VDDHD VDDI PCH L=60N W=1U M=1
MM14 LWDT[1] GWDT_YL VDDHD VDDI PCH L=60N W=1U M=1
MM24 GWDC_YL YL[1] VDDHD VDDI PCH L=60N W=300N M=1
MM13 GWDT_YL GW VDDHD VDDI PCH L=60N W=300N M=1
MM6 SAE_OFF SAE_OFFB VDDHD VDDI PCH L=60N W=300N M=1
MM19 GWDT_YLB GW VDDHD VDDI PCH L=60N W=300N M=1
MM12 GWDT_YL YL[1] VDDHD VDDI PCH L=60N W=300N M=1
MM32 GWDC_YLB YL[0] VDDHD VDDI PCH L=60N W=300N M=1
MM20 GWDT_YLB YL[0] VDDHD VDDI PCH L=60N W=300N M=1
MM18 LWDT[0] GWDT_YLB VDDHD VDDI PCH L=60N W=1U M=1
MM38 WC[0] LWDT[0] VDDHD VDDI PCH L=65.0N W=500N M=4
MM37 WT[1] LWDC[1] VDDHD VDDI PCH L=65.0N W=500N M=4
MM1 WT[0] LWDC[0] VDDHD VDDI PCH L=65.0N W=500N M=4
MM10 SAE_OFFB GBLB VDDHD VDDI PCH L=60N W=300N M=1
MM11 SAE_OFFB GBL VDDHD VDDI PCH L=60N W=300N M=1
MM40 WC[1] LWDT[1] VDDHD VDDI PCH L=65.0N W=500N M=4
MM41 WC[1] LWDT[1] VSSI VSSI NCH L=65.0N W=1.5U M=4
MM27 NET0588 YL[1] VSSI VSSI NCH L=60N W=300N M=1
MM28 GWDC_YL GWB NET0588 VSSI NCH L=60N W=300N M=1
MM29 LWDC[1] GWDC_YL VSSI VSSI NCH L=60N W=500N M=1
MM35 NET0568 YL[0] VSSI VSSI NCH L=60N W=300N M=1
MM15 NET0290 YL[1] VSSI VSSI NCH L=60N W=300N M=1
MM16 GWDT_YL GW NET0290 VSSI NCH L=60N W=300N M=1
MM23 NET0270 YL[0] VSSI VSSI NCH L=60N W=300N M=1
MM22 GWDT_YLB GW NET0270 VSSI NCH L=60N W=300N M=1
MM7 SAE_OFF SAE_OFFB VSSI VSSI NCH L=60N W=300N M=1
MM8 SAE_OFFB GBL NET244 VSSI NCH L=60N W=300N M=1
MM9 NET244 GBLB VSSI VSSI NCH L=60N W=300N M=1
MM17 LWDT[1] GWDT_YL VSSI VSSI NCH L=60N W=500N M=1
MM33 LWDC[0] GWDC_YLB VSSI VSSI NCH L=60N W=500N M=1
MM34 GWDC_YLB GWB NET0568 VSSI NCH L=60N W=300N M=1
MM36 WT[1] LWDC[1] VSSI VSSI NCH L=65.0N W=1.5U M=4
MM21 LWDT[0] GWDT_YLB VSSI VSSI NCH L=60N W=500N M=1
MM39 WC[0] LWDT[0] VSSI VSSI NCH L=65.0N W=1.5U M=4
MM0 WT[0] LWDC[0] VSSI VSSI NCH L=65.0N W=1.5U M=4
XI248 SAEC VSSI VDDI SAE S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.6U LP=0.06U M=1
XI105 RE VSSI VDDI WRITE S1AHSF400W40_AINV FN=3 WN=0.5U LN=0.07U FP=3 WP=1U LP=0.07U M=1
XINV4 WE VSSI VDDI READ S1AHSF400W40_AINV FN=3 WN=0.5U LN=0.07U FP=3 WP=1U LP=0.07U M=1
XI235 SAEB SAE_OFF VSSI VDDI SAEC S1AHSF400W40_ANAND FN2=1 WN2=0.25U LN2=0.06U FN1=1 
+ WN1=0.25U LN1=0.06U FP1=1 WP1=0.25U LP1=0.06U FP2=1 WP2=0.25U LP2=0.06U M=1
XI75 BLEQB_UP_0 YL[0] VSSI VDDI PGB_UP_0 S1AHSF400W40_ANAND FN2=1 WN2=0.5U LN2=0.06U 
+ FN1=1 WN1=0.5U LN1=0.06U FP1=1 WP1=0.5U LP1=0.06U FP2=1 WP2=0.5U LP2=0.06U 
+ M=1
XI77 BLEQB_DN_0 YL[0] VSSI VDDI PGB_DN_0 S1AHSF400W40_ANAND FN2=1 WN2=0.5U LN2=0.06U 
+ FN1=1 WN1=0.5U LN1=0.06U FP1=1 WP1=0.5U LP1=0.06U FP2=1 WP2=0.5U LP2=0.06U 
+ M=1
XI78 BLEQB_DN_1 YL[1] VSSI VDDI PGB_DN_1 S1AHSF400W40_ANAND FN2=1 WN2=0.5U LN2=0.06U 
+ FN1=1 WN1=0.5U LN1=0.06U FP1=1 WP1=0.5U LP1=0.06U FP2=1 WP2=0.5U LP2=0.06U 
+ M=1
XI76 BLEQB_UP_1 YL[1] VSSI VDDI PGB_UP_1 S1AHSF400W40_ANAND FN2=1 WN2=0.5U LN2=0.06U 
+ FN1=1 WN1=0.5U LN1=0.06U FP1=1 WP1=0.5U LP1=0.06U FP2=1 WP2=0.5U LP2=0.06U 
+ M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LIO_M16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LIO_M16 BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_DN[4] BLB_DN[5] 
+ BLB_DN[6] BLB_DN[7] BLB_DN[8] BLB_DN[9] BLB_DN[10] BLB_DN[11] BLB_DN[12] 
+ BLB_DN[13] BLB_DN[14] BLB_DN[15] BLB_UP[0] BLB_UP[1] BLB_UP[2] BLB_UP[3] 
+ BLB_UP[4] BLB_UP[5] BLB_UP[6] BLB_UP[7] BLB_UP[8] BLB_UP[9] BLB_UP[10] 
+ BLB_UP[11] BLB_UP[12] BLB_UP[13] BLB_UP[14] BLB_UP[15] BLEQ_DN BLEQ_UP 
+ BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] BL_DN[4] BL_DN[5] BL_DN[6] BL_DN[7] 
+ BL_DN[8] BL_DN[9] BL_DN[10] BL_DN[11] BL_DN[12] BL_DN[13] BL_DN[14] 
+ BL_DN[15] BL_UP[0] BL_UP[1] BL_UP[2] BL_UP[3] BL_UP[4] BL_UP[5] BL_UP[6] 
+ BL_UP[7] BL_UP[8] BL_UP[9] BL_UP[10] BL_UP[11] BL_UP[12] BL_UP[13] BL_UP[14] 
+ BL_UP[15] GBL GBLB GW GWB RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] 
+ Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] 
+ Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
*.PININFO BLEQ_DN:I BLEQ_UP:I GW:I GWB:I RE:I SAEB:I WE:I YL_LIO[0]:I 
*.PININFO YL_LIO[1]:I Y_DN[0]:I Y_DN[1]:I Y_DN[2]:I Y_DN[3]:I Y_DN[4]:I 
*.PININFO Y_DN[5]:I Y_DN[6]:I Y_DN[7]:I Y_UP[0]:I Y_UP[1]:I Y_UP[2]:I 
*.PININFO Y_UP[3]:I Y_UP[4]:I Y_UP[5]:I Y_UP[6]:I Y_UP[7]:I BLB_DN[0]:B 
*.PININFO BLB_DN[1]:B BLB_DN[2]:B BLB_DN[3]:B BLB_DN[4]:B BLB_DN[5]:B 
*.PININFO BLB_DN[6]:B BLB_DN[7]:B BLB_DN[8]:B BLB_DN[9]:B BLB_DN[10]:B 
*.PININFO BLB_DN[11]:B BLB_DN[12]:B BLB_DN[13]:B BLB_DN[14]:B BLB_DN[15]:B 
*.PININFO BLB_UP[0]:B BLB_UP[1]:B BLB_UP[2]:B BLB_UP[3]:B BLB_UP[4]:B 
*.PININFO BLB_UP[5]:B BLB_UP[6]:B BLB_UP[7]:B BLB_UP[8]:B BLB_UP[9]:B 
*.PININFO BLB_UP[10]:B BLB_UP[11]:B BLB_UP[12]:B BLB_UP[13]:B BLB_UP[14]:B 
*.PININFO BLB_UP[15]:B BL_DN[0]:B BL_DN[1]:B BL_DN[2]:B BL_DN[3]:B BL_DN[4]:B 
*.PININFO BL_DN[5]:B BL_DN[6]:B BL_DN[7]:B BL_DN[8]:B BL_DN[9]:B BL_DN[10]:B 
*.PININFO BL_DN[11]:B BL_DN[12]:B BL_DN[13]:B BL_DN[14]:B BL_DN[15]:B 
*.PININFO BL_UP[0]:B BL_UP[1]:B BL_UP[2]:B BL_UP[3]:B BL_UP[4]:B BL_UP[5]:B 
*.PININFO BL_UP[6]:B BL_UP[7]:B BL_UP[8]:B BL_UP[9]:B BL_UP[10]:B BL_UP[11]:B 
*.PININFO BL_UP[12]:B BL_UP[13]:B BL_UP[14]:B BL_UP[15]:B GBL:B GBLB:B VDDHD:B 
*.PININFO VDDI:B VSSI:B
XYPASS_DN_1 BL_DN[8] BL_DN[9] BL_DN[10] BL_DN[11] BL_DN[12] BL_DN[13] 
+ BL_DN[14] BL_DN[15] BLB_DN[8] BLB_DN[9] BLB_DN[10] BLB_DN[11] BLB_DN[12] 
+ BLB_DN[13] BLB_DN[14] BLB_DN[15] BLEQ_DN BLEQB_DN_1 DL_DN_1 DLB_DN_1 READ 
+ VDDI VSSI WC[1] WRITE WT[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] 
+ Y_DN[6] Y_DN[7] S1AHSF400W40_YPASS_M8
XYPASS_DN_0 BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] BL_DN[4] BL_DN[5] BL_DN[6] 
+ BL_DN[7] BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_DN[4] BLB_DN[5] 
+ BLB_DN[6] BLB_DN[7] BLEQ_DN BLEQB_DN_0 DL_DN_0 DLB_DN_0 READ VDDI VSSI WC[0] 
+ WRITE WT[0] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] 
+ S1AHSF400W40_YPASS_M8
XYPASS_UP_0 BL_UP[0] BL_UP[1] BL_UP[2] BL_UP[3] BL_UP[4] BL_UP[5] BL_UP[6] 
+ BL_UP[7] BLB_UP[0] BLB_UP[1] BLB_UP[2] BLB_UP[3] BLB_UP[4] BLB_UP[5] 
+ BLB_UP[6] BLB_UP[7] BLEQ_UP BLEQB_UP_0 DL_UP_0 DLB_UP_0 READ VDDI VSSI WC[0] 
+ WRITE WT[0] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] 
+ S1AHSF400W40_YPASS_M8
XYPASS_UP_1 BL_UP[8] BL_UP[9] BL_UP[10] BL_UP[11] BL_UP[12] BL_UP[13] 
+ BL_UP[14] BL_UP[15] BLB_UP[8] BLB_UP[9] BLB_UP[10] BLB_UP[11] BLB_UP[12] 
+ BLB_UP[13] BLB_UP[14] BLB_UP[15] BLEQ_UP BLEQB_UP_1 DL_UP_1 DLB_UP_1 READ 
+ VDDI VSSI WC[1] WRITE WT[1] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] 
+ Y_UP[6] Y_UP[7] S1AHSF400W40_YPASS_M8
XIO_RWBLK BLEQB_DN_0 BLEQB_DN_1 BLEQB_UP_0 BLEQB_UP_1 BLEQ_DN BLEQ_UP DLB_DN_0 
+ DLB_DN_1 DLB_UP_0 DLB_UP_1 DL_DN_0 DL_DN_1 DL_UP_0 DL_UP_1 GBL GBLB GW GWB 
+ RE READ SAEB VDDHD VDDI VSSI WC[0] WC[1] WE WRITE WT[0] WT[1] YL_LIO[0] 
+ YL_LIO[1] S1AHSF400W40_IO_RWBLK_M16
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    SA_M8
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SA_M8 DLB_DN DLB_UP DL_DN DL_UP GBL GBLB PGB_DN PGB_UP PREB SAE VDDI 
+ VSSI
*.PININFO PGB_DN:I PGB_UP:I PREB:I SAE:I DLB_DN:B DLB_UP:B DL_DN:B DL_UP:B 
*.PININFO GBL:B GBLB:B VDDI:B VSSI:B
MP11 DLB_IN PREB VDDI VDDI PCH L=100N W=1U M=1
MP7 DLB_IN PGB_UP DLB_UP VDDI PCH L=100N W=1U M=1
MP8 DL_IN PREB DLB_IN VDDI PCH L=120.0N W=1U M=2
MP3 DLB_IN DL_IN VDDI VDDI PCH L=120.0N W=1U M=1
MP14 DLB_IN PGB_DN DLB_DN VDDI PCH L=100N W=1U M=1
MP2 VDDI DLB_IN DL_IN VDDI PCH L=120.0N W=1U M=1
MP13 DL_DN PGB_DN DL_IN VDDI PCH L=100N W=1U M=1
MP6 DL_UP PGB_UP DL_IN VDDI PCH L=100N W=1U M=1
MP10 DL_IN PREB VDDI VDDI PCH L=100N W=1U M=1
MN12 GBLB SOB VSSI VSSI NCH L=65.0N W=2.5U M=2
MN11 GBL SO VSSI VSSI NCH L=65.0N W=2.5U M=2
MN1 DLB_IN DL_IN NS VSSI NCH L=180.0N W=500N M=4
MN0 NS DLB_IN DL_IN VSSI NCH L=180.0N W=500N M=4
MN2 NS SAE VSSI VSSI NCH L=80N W=500N M=4
XINV0 DL_IN VSSI VDDI SO S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U LP=0.06U M=1
XINV1 DLB_IN VSSI VDDI SOB S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    IO_RWBLK_M8
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_IO_RWBLK_M8 BLEQB_DN BLEQB_UP BLEQ_DN BLEQ_UP DLB_DN DLB_UP DL_DN 
+ DL_UP GBL GBLB GW GWB RE READ SAEB VDDHD VDDI VSSI WC WE WRITE WT
*.PININFO BLEQB_DN:I BLEQB_UP:I BLEQ_DN:I BLEQ_UP:I GW:I GWB:I RE:I SAEB:I 
*.PININFO WE:I READ:O WC:O WRITE:O WT:O DLB_DN:B DLB_UP:B DL_DN:B DL_UP:B 
*.PININFO GBL:B GBLB:B VDDHD:B VDDI:B VSSI:B
XI235 SAEB SAE_OFF VSSI VDDI SAEC S1AHSF400W40_ANAND FN2=1 WN2=0.25U LN2=0.06U FN1=1 
+ WN1=0.25U LN1=0.06U FP1=1 WP1=0.25U LP1=0.06U FP2=1 WP2=0.25U LP2=0.06U M=1
XI222 SAEC BLEQ_UP BLEQ_DN VSSI VDDI PREB S1AHSF400W40_ANAND3 FN3=1 WN3=0.4U LN3=0.06U 
+ FN2=1 WN2=0.4U LN2=0.06U FN1=1 WN1=0.4U LN1=0.06U FP1=1 WP1=0.4U LP1=0.06U 
+ FP2=1 WP2=0.4U LP2=0.06U FP3=1 WP3=0.4U LP3=0.06U M=1
MM3 WC GW VDDHD VDDI PCH L=65.0N W=500N M=4
MM6 SAE_OFF SAE_OFFB VDDHD VDDI PCH L=60N W=300N M=1
MM10 SAE_OFFB GBLB VDDHD VDDI PCH L=60N W=300N M=1
MM11 SAE_OFFB GBL VDDHD VDDI PCH L=60N W=300N M=1
MM1 WT GWB VDDHD VDDI PCH L=65.0N W=500N M=4
MM2 WC GW VSSI VSSI NCH L=65.0N W=1.5U M=4
MM9 NET150 GBLB VSSI VSSI NCH L=60N W=300N M=1
MM7 SAE_OFF SAE_OFFB VSSI VSSI NCH L=60N W=300N M=1
MM8 SAE_OFFB GBL NET150 VSSI NCH L=60N W=300N M=1
MM0 WT GWB VSSI VSSI NCH L=65.0N W=1.5U M=4
XI248 SAEC VSSI VDDI SAE S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.6U LP=0.06U M=1
XI273 BLEQB_DN VSSI VDDI PGB_DN S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=0.36U 
+ LP=0.06U M=1
XI272 BLEQB_UP VSSI VDDI PGB_UP S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=0.36U 
+ LP=0.06U M=1
XI234 RE VSSI VDDI WRITE S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.07U FP=1 WP=1U LP=0.07U M=1
XI268 WE VSSI VDDI READ S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.07U FP=1 WP=1U LP=0.07U M=1
XSA DLB_DN DLB_UP DL_DN DL_UP GBL GBLB PGB_DN PGB_UP PREB SAE VDDI VSSI S1AHSF400W40_SA_M8
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LIO_M8
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LIO_M8 BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_DN[4] BLB_DN[5] 
+ BLB_DN[6] BLB_DN[7] BLB_UP[0] BLB_UP[1] BLB_UP[2] BLB_UP[3] BLB_UP[4] 
+ BLB_UP[5] BLB_UP[6] BLB_UP[7] BLEQ_DN BLEQ_UP BL_DN[0] BL_DN[1] BL_DN[2] 
+ BL_DN[3] BL_DN[4] BL_DN[5] BL_DN[6] BL_DN[7] BL_UP[0] BL_UP[1] BL_UP[2] 
+ BL_UP[3] BL_UP[4] BL_UP[5] BL_UP[6] BL_UP[7] GBL GBLB GW GWB RE SAEB VDDHD 
+ VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] 
+ Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] 
+ Y_UP[6] Y_UP[7]
*.PININFO BLEQ_DN:I BLEQ_UP:I GW:I GWB:I RE:I SAEB:I WE:I YL_LIO[0]:I 
*.PININFO YL_LIO[1]:I Y_DN[0]:I Y_DN[1]:I Y_DN[2]:I Y_DN[3]:I Y_DN[4]:I 
*.PININFO Y_DN[5]:I Y_DN[6]:I Y_DN[7]:I Y_UP[0]:I Y_UP[1]:I Y_UP[2]:I 
*.PININFO Y_UP[3]:I Y_UP[4]:I Y_UP[5]:I Y_UP[6]:I Y_UP[7]:I BLB_DN[0]:B 
*.PININFO BLB_DN[1]:B BLB_DN[2]:B BLB_DN[3]:B BLB_DN[4]:B BLB_DN[5]:B 
*.PININFO BLB_DN[6]:B BLB_DN[7]:B BLB_UP[0]:B BLB_UP[1]:B BLB_UP[2]:B 
*.PININFO BLB_UP[3]:B BLB_UP[4]:B BLB_UP[5]:B BLB_UP[6]:B BLB_UP[7]:B 
*.PININFO BL_DN[0]:B BL_DN[1]:B BL_DN[2]:B BL_DN[3]:B BL_DN[4]:B BL_DN[5]:B 
*.PININFO BL_DN[6]:B BL_DN[7]:B BL_UP[0]:B BL_UP[1]:B BL_UP[2]:B BL_UP[3]:B 
*.PININFO BL_UP[4]:B BL_UP[5]:B BL_UP[6]:B BL_UP[7]:B GBL:B GBLB:B VDDHD:B 
*.PININFO VDDI:B VSSI:B
XIO_RWBLK BLEQB_DN_0 BLEQB_UP_0 BLEQ_DN BLEQ_UP DLB_DN DLB_UP DL_DN DL_UP GBL 
+ GBLB GW GWB RE READ SAEB VDDHD VDDI VSSI WC WE WRITE WT S1AHSF400W40_IO_RWBLK_M8
XYPASS_DN BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] BL_DN[4] BL_DN[5] BL_DN[6] 
+ BL_DN[7] BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_DN[4] BLB_DN[5] 
+ BLB_DN[6] BLB_DN[7] BLEQ_DN BLEQB_DN_0 DL_DN DLB_DN READ VDDI VSSI WC WRITE 
+ WT Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] S1AHSF400W40_YPASS_M8
XYPASS_UP BL_UP[0] BL_UP[1] BL_UP[2] BL_UP[3] BL_UP[4] BL_UP[5] BL_UP[6] 
+ BL_UP[7] BLB_UP[0] BLB_UP[1] BLB_UP[2] BLB_UP[3] BLB_UP[4] BLB_UP[5] 
+ BLB_UP[6] BLB_UP[7] BLEQ_UP BLEQB_UP_0 DL_UP DLB_UP READ VDDI VSSI WC WRITE 
+ WT Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_YPASS_M8
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    SA_M4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SA_M4 DLB_DN DLB_UP DL_DN DL_UP GBL GBLB PGB_DN PGB_UP PREB SAE VDDI 
+ VSSI
*.PININFO PGB_DN:I PGB_UP:I PREB:I SAE:I DLB_DN:B DLB_UP:B DL_DN:B DL_UP:B 
*.PININFO GBL:B GBLB:B VDDI:B VSSI:B
MP11 DLB_IN PREB VDDI VDDI PCH L=100N W=1U M=1
MP8 DL_IN PREB DLB_IN VDDI PCH L=120.0N W=1U M=2
MP3 DLB_IN DL_IN VDDI VDDI PCH L=120.0N W=1U M=1
MP13 DL_DN PGB_DN DL_IN VDDI PCH L=100N W=1U M=1
MP2 VDDI DLB_IN DL_IN VDDI PCH L=120.0N W=1U M=1
MP7 DLB_IN PGB_UP DLB_UP VDDI PCH L=100N W=1U M=1
MP14 DLB_IN PGB_DN DLB_DN VDDI PCH L=100N W=1U M=1
MP6 DL_UP PGB_UP DL_IN VDDI PCH L=100N W=1U M=1
MP10 DL_IN PREB VDDI VDDI PCH L=100N W=1U M=1
MN12 GBLB SOB VSSI VSSI NCH L=60N W=600N M=8
MN11 GBL SO VSSI VSSI NCH L=60N W=600N M=8
MN0 NS DLB_IN DL_IN VSSI NCH L=180.0N W=500N M=4
MN1 DLB_IN DL_IN NS VSSI NCH L=180.0N W=500N M=4
MN2 NS SAE VSSI VSSI NCH L=80N W=500N M=4
XINV0 DL_IN VSSI VDDI SO S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U LP=0.06U M=1
XINV1 DLB_IN VSSI VDDI SOB S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    IO_RWBLK_M4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_IO_RWBLK_M4 BLEQB_DN BLEQB_UP BLEQ_DN BLEQ_UP DLB_DN DLB_UP DL_DN 
+ DL_UP GBL GBLB GW GWB SAEB VDDHD VDDI VSSI WC WT
*.PININFO BLEQB_DN:I BLEQB_UP:I BLEQ_DN:I BLEQ_UP:I GW:I GWB:I SAEB:I WC:O 
*.PININFO WT:O DLB_DN:B DLB_UP:B DL_DN:B DL_UP:B GBL:B GBLB:B VDDHD:B VDDI:B 
*.PININFO VSSI:B
XSA DLB_DN DLB_UP DL_DN DL_UP GBL GBLB PGB_DN PGB_UP PREB SAE VDDI VSSI S1AHSF400W40_SA_M4
XI222 SAEC BLEQ_UP BLEQ_DN VSSI VDDI PREB S1AHSF400W40_ANAND3 FN3=1 WN3=0.4U LN3=0.06U 
+ FN2=1 WN2=0.4U LN2=0.06U FN1=1 WN1=0.4U LN1=0.06U FP1=1 WP1=0.4U LP1=0.06U 
+ FP2=1 WP2=0.4U LP2=0.06U FP3=1 WP3=0.4U LP3=0.06U M=1
MM6 SAE_OFF SAE_OFFB VDDHD VDDI PCH L=60N W=300N M=2
MM10 SAE_OFFB GBLB VDDHD VDDI PCH L=60N W=300N M=1
MM11 SAE_OFFB GBL VDDHD VDDI PCH L=60N W=300N M=1
MP27 WC GW VDDHD VDDI PCH L=60N W=330.0N M=5
MP25 WT GWB VDDHD VDDI PCH L=60N W=330.0N M=5
MM9 NET117 GBLB VSSI VSSI NCH L=60N W=300N M=1
MM7 SAE_OFF SAE_OFFB VSSI VSSI NCH L=60N W=300N M=1
MM8 SAE_OFFB GBL NET117 VSSI NCH L=60N W=300N M=1
MN13 WT GWB VSSI VSSI NCH L=60N W=990.0N M=5
MN0 WC GW VSSI VSSI NCH L=60N W=990.0N M=5
XI235 SAEB SAE_OFF VSSI VDDI SAEC S1AHSF400W40_ANAND FN2=1 WN2=0.25U LN2=0.06U FN1=1 
+ WN1=0.25U LN1=0.06U FP1=1 WP1=0.25U LP1=0.06U FP2=1 WP2=0.25U LP2=0.06U M=1
XI54 BLEQB_DN VSSI VDDI PGB_DN S1AHSF400W40_AINV FN=1 WN=0.36U LN=0.06U FP=1 WP=0.36U 
+ LP=0.06U M=1
XI58 BLEQB_UP VSSI VDDI PGB_UP S1AHSF400W40_AINV FN=1 WN=0.36U LN=0.06U FP=1 WP=0.36U 
+ LP=0.06U M=1
XI248 SAEC VSSI VDDI SAE S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.6U LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    YPASS_M4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_YPASS_M4 BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] BLEQ 
+ BLEQB DL DLB VDDI VSSI WC WT Y[0] Y[1] Y[2] Y[3] Y[4] Y[5] Y[6] Y[7]
*.PININFO BLEQ:I Y[0]:I Y[1]:I Y[2]:I Y[3]:I Y[4]:I Y[5]:I Y[6]:I Y[7]:I 
*.PININFO BL[0]:B BL[1]:B BL[2]:B BL[3]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B 
*.PININFO BLEQB:B DL:B DLB:B VDDI:B VSSI:B WC:B WT:B
XI284<0> BLB[0] BL[0] BLEQB VDDI S1AHSF400W40_PRECHARGE
XI284<1> BLB[1] BL[1] BLEQB VDDI S1AHSF400W40_PRECHARGE
XI284<2> BLB[2] BL[2] BLEQB VDDI S1AHSF400W40_PRECHARGE
XI284<3> BLB[3] BL[3] BLEQB VDDI S1AHSF400W40_PRECHARGE
MP22 VDDI BLEQB DL VDDI PCH L=60N W=200N M=1
MM2<0> DL YB[0] BL[0] VDDI PCH L=60N W=800N M=1
MM2<1> DL YB[1] BL[1] VDDI PCH L=60N W=800N M=1
MM2<2> DL YB[2] BL[2] VDDI PCH L=60N W=800N M=1
MM2<3> DL YB[3] BL[3] VDDI PCH L=60N W=800N M=1
MP3 DLB BLEQB VDDI VDDI PCH L=60N W=200N M=1
MM3<0> DLB YB[0] BLB[0] VDDI PCH L=60N W=800N M=1
MM3<1> DLB YB[1] BLB[1] VDDI PCH L=60N W=800N M=1
MM3<2> DLB YB[2] BLB[2] VDDI PCH L=60N W=800N M=1
MM3<3> DLB YB[3] BLB[3] VDDI PCH L=60N W=800N M=1
MN18<0> BLB[0] Y[4] WC VSSI NCH L=60N W=1.6U M=1
MN18<1> BLB[1] Y[5] WC VSSI NCH L=60N W=1.6U M=1
MN18<2> BLB[2] Y[6] WC VSSI NCH L=60N W=1.6U M=1
MN18<3> BLB[3] Y[7] WC VSSI NCH L=60N W=1.6U M=1
MM4<0> BL[0] Y[4] WT VSSI NCH L=60N W=1.6U M=1
MM4<1> BL[1] Y[5] WT VSSI NCH L=60N W=1.6U M=1
MM4<2> BL[2] Y[6] WT VSSI NCH L=60N W=1.6U M=1
MM4<3> BL[3] Y[7] WT VSSI NCH L=60N W=1.6U M=1
XI285 BLEQ VSSI VDDI BLEQB S1AHSF400W40_AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=1.6U LP=0.06U 
+ M=1
XND0<0> Y[0] VSSI VDDI YB[0] S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.3U 
+ LP=0.06U M=1
XND0<1> Y[1] VSSI VDDI YB[1] S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.3U 
+ LP=0.06U M=1
XND0<2> Y[2] VSSI VDDI YB[2] S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.3U 
+ LP=0.06U M=1
XND0<3> Y[3] VSSI VDDI YB[3] S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.3U 
+ LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LIO_M4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LIO_M4 BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_UP[0] BLB_UP[1] 
+ BLB_UP[2] BLB_UP[3] BLEQ_DN BLEQ_UP BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] 
+ BL_UP[0] BL_UP[1] BL_UP[2] BL_UP[3] GBL GBLB GW GWB RE SAEB VDDHD VDDI VSSI 
+ WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] 
+ Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] 
+ Y_UP[7]
*.PININFO BLEQ_DN:I BLEQ_UP:I GW:I GWB:I RE:I SAEB:I WE:I YL_LIO[0]:I 
*.PININFO YL_LIO[1]:I Y_DN[0]:I Y_DN[1]:I Y_DN[2]:I Y_DN[3]:I Y_DN[4]:I 
*.PININFO Y_DN[5]:I Y_DN[6]:I Y_DN[7]:I Y_UP[0]:I Y_UP[1]:I Y_UP[2]:I 
*.PININFO Y_UP[3]:I Y_UP[4]:I Y_UP[5]:I Y_UP[6]:I Y_UP[7]:I BLB_DN[0]:B 
*.PININFO BLB_DN[1]:B BLB_DN[2]:B BLB_DN[3]:B BLB_UP[0]:B BLB_UP[1]:B 
*.PININFO BLB_UP[2]:B BLB_UP[3]:B BL_DN[0]:B BL_DN[1]:B BL_DN[2]:B BL_DN[3]:B 
*.PININFO BL_UP[0]:B BL_UP[1]:B BL_UP[2]:B BL_UP[3]:B GBL:B GBLB:B VDDHD:B 
*.PININFO VDDI:B VSSI:B
XIO_RWBLK BLEQB_DN_0 BLEQB_UP_0 BLEQ_DN BLEQ_UP DLB_DN DLB_UP DL_DN DL_UP GBL 
+ GBLB GW GWB SAEB VDDHD VDDI VSSI WC WT S1AHSF400W40_IO_RWBLK_M4
XYPASS_D BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] BLB_DN[0] BLB_DN[1] BLB_DN[2] 
+ BLB_DN[3] BLEQ_DN BLEQB_DN_0 DL_DN DLB_DN VDDI VSSI WC WT Y_DN[0] Y_DN[1] 
+ Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] S1AHSF400W40_YPASS_M4
XYPASS_U BL_UP[0] BL_UP[1] BL_UP[2] BL_UP[3] BLB_UP[0] BLB_UP[1] BLB_UP[2] 
+ BLB_UP[3] BLEQ_UP BLEQB_UP_0 DL_UP DLB_UP VDDI VSSI WC WT Y_UP[0] Y_UP[1] 
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_YPASS_M4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    ARR_LIO_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ARR_LIO_SIM BLB_DN_BT[0] BLB_DN_BT[1] BLB_DN_BT[2] BLB_DN_BT[3] 
+ BLB_DN_BT[4] BLB_DN_BT[5] BLB_DN_BT[6] BLB_DN_BT[7] BLB_DN_BT[8] 
+ BLB_DN_BT[9] BLB_DN_BT[10] BLB_DN_BT[11] BLB_DN_BT[12] BLB_DN_BT[13] 
+ BLB_DN_BT[14] BLB_DN_BT[15] BLB_UP_TP[0] BLB_UP_TP[1] BLB_UP_TP[2] 
+ BLB_UP_TP[3] BLB_UP_TP[4] BLB_UP_TP[5] BLB_UP_TP[6] BLB_UP_TP[7] 
+ BLB_UP_TP[8] BLB_UP_TP[9] BLB_UP_TP[10] BLB_UP_TP[11] BLB_UP_TP[12] 
+ BLB_UP_TP[13] BLB_UP_TP[14] BLB_UP_TP[15] BLEQ_DN_LT BLEQ_DN_RT BLEQ_UP_LT 
+ BLEQ_UP_RT BL_DN_BT[0] BL_DN_BT[1] BL_DN_BT[2] BL_DN_BT[3] BL_DN_BT[4] 
+ BL_DN_BT[5] BL_DN_BT[6] BL_DN_BT[7] BL_DN_BT[8] BL_DN_BT[9] BL_DN_BT[10] 
+ BL_DN_BT[11] BL_DN_BT[12] BL_DN_BT[13] BL_DN_BT[14] BL_DN_BT[15] BL_UP_TP[0] 
+ BL_UP_TP[1] BL_UP_TP[2] BL_UP_TP[3] BL_UP_TP[4] BL_UP_TP[5] BL_UP_TP[6] 
+ BL_UP_TP[7] BL_UP_TP[8] BL_UP_TP[9] BL_UP_TP[10] BL_UP_TP[11] BL_UP_TP[12] 
+ BL_UP_TP[13] BL_UP_TP[14] BL_UP_TP[15] CVDDI GBLB_BT GBLB_TP GBL_BT GBL_TP 
+ GWB_BT GWB_TP GW_BT GW_TP RE_LT RE_RT SAEB_LT SAEB_RT VDDHD VDDI VSSI WE_LT 
+ WE_RT YL_LIO_LT[0] YL_LIO_LT[1] YL_LIO_RT[0] YL_LIO_RT[1] Y_DN_LT[0] 
+ Y_DN_LT[1] Y_DN_LT[2] Y_DN_LT[3] Y_DN_LT[4] Y_DN_LT[5] Y_DN_LT[6] Y_DN_LT[7] 
+ Y_DN_RT[0] Y_DN_RT[1] Y_DN_RT[2] Y_DN_RT[3] Y_DN_RT[4] Y_DN_RT[5] Y_DN_RT[6] 
+ Y_DN_RT[7] Y_UP_LT[0] Y_UP_LT[1] Y_UP_LT[2] Y_UP_LT[3] Y_UP_LT[4] Y_UP_LT[5] 
+ Y_UP_LT[6] Y_UP_LT[7] Y_UP_RT[0] Y_UP_RT[1] Y_UP_RT[2] Y_UP_RT[3] Y_UP_RT[4] 
+ Y_UP_RT[5] Y_UP_RT[6] Y_UP_RT[7]
*.PININFO BLB_DN_BT[0]:B BLB_DN_BT[1]:B BLB_DN_BT[2]:B BLB_DN_BT[3]:B 
*.PININFO BLB_DN_BT[4]:B BLB_DN_BT[5]:B BLB_DN_BT[6]:B BLB_DN_BT[7]:B 
*.PININFO BLB_DN_BT[8]:B BLB_DN_BT[9]:B BLB_DN_BT[10]:B BLB_DN_BT[11]:B 
*.PININFO BLB_DN_BT[12]:B BLB_DN_BT[13]:B BLB_DN_BT[14]:B BLB_DN_BT[15]:B 
*.PININFO BLB_UP_TP[0]:B BLB_UP_TP[1]:B BLB_UP_TP[2]:B BLB_UP_TP[3]:B 
*.PININFO BLB_UP_TP[4]:B BLB_UP_TP[5]:B BLB_UP_TP[6]:B BLB_UP_TP[7]:B 
*.PININFO BLB_UP_TP[8]:B BLB_UP_TP[9]:B BLB_UP_TP[10]:B BLB_UP_TP[11]:B 
*.PININFO BLB_UP_TP[12]:B BLB_UP_TP[13]:B BLB_UP_TP[14]:B BLB_UP_TP[15]:B 
*.PININFO BLEQ_DN_LT:B BLEQ_DN_RT:B BLEQ_UP_LT:B BLEQ_UP_RT:B BL_DN_BT[0]:B 
*.PININFO BL_DN_BT[1]:B BL_DN_BT[2]:B BL_DN_BT[3]:B BL_DN_BT[4]:B 
*.PININFO BL_DN_BT[5]:B BL_DN_BT[6]:B BL_DN_BT[7]:B BL_DN_BT[8]:B 
*.PININFO BL_DN_BT[9]:B BL_DN_BT[10]:B BL_DN_BT[11]:B BL_DN_BT[12]:B 
*.PININFO BL_DN_BT[13]:B BL_DN_BT[14]:B BL_DN_BT[15]:B BL_UP_TP[0]:B 
*.PININFO BL_UP_TP[1]:B BL_UP_TP[2]:B BL_UP_TP[3]:B BL_UP_TP[4]:B 
*.PININFO BL_UP_TP[5]:B BL_UP_TP[6]:B BL_UP_TP[7]:B BL_UP_TP[8]:B 
*.PININFO BL_UP_TP[9]:B BL_UP_TP[10]:B BL_UP_TP[11]:B BL_UP_TP[12]:B 
*.PININFO BL_UP_TP[13]:B BL_UP_TP[14]:B BL_UP_TP[15]:B CVDDI:B GBLB_BT:B 
*.PININFO GBLB_TP:B GBL_BT:B GBL_TP:B GWB_BT:B GWB_TP:B GW_BT:B GW_TP:B 
*.PININFO RE_LT:B RE_RT:B SAEB_LT:B SAEB_RT:B VDDHD:B VDDI:B VSSI:B WE_LT:B 
*.PININFO WE_RT:B YL_LIO_LT[0]:B YL_LIO_LT[1]:B YL_LIO_RT[0]:B YL_LIO_RT[1]:B 
*.PININFO Y_DN_LT[0]:B Y_DN_LT[1]:B Y_DN_LT[2]:B Y_DN_LT[3]:B Y_DN_LT[4]:B 
*.PININFO Y_DN_LT[5]:B Y_DN_LT[6]:B Y_DN_LT[7]:B Y_DN_RT[0]:B Y_DN_RT[1]:B 
*.PININFO Y_DN_RT[2]:B Y_DN_RT[3]:B Y_DN_RT[4]:B Y_DN_RT[5]:B Y_DN_RT[6]:B 
*.PININFO Y_DN_RT[7]:B Y_UP_LT[0]:B Y_UP_LT[1]:B Y_UP_LT[2]:B Y_UP_LT[3]:B 
*.PININFO Y_UP_LT[4]:B Y_UP_LT[5]:B Y_UP_LT[6]:B Y_UP_LT[7]:B Y_UP_RT[0]:B 
*.PININFO Y_UP_RT[1]:B Y_UP_RT[2]:B Y_UP_RT[3]:B Y_UP_RT[4]:B Y_UP_RT[5]:B 
*.PININFO Y_UP_RT[6]:B Y_UP_RT[7]:B
XLIO_M16 NET040[0] NET040[1] NET040[2] NET040[3] NET040[4] NET040[5] NET040[6] 
+ NET040[7] NET040[8] NET040[9] NET040[10] NET040[11] NET040[12] NET040[13] 
+ NET040[14] NET040[15] NET038[0] NET038[1] NET038[2] NET038[3] NET038[4] 
+ NET038[5] NET038[6] NET038[7] NET038[8] NET038[9] NET038[10] NET038[11] 
+ NET038[12] NET038[13] NET038[14] NET038[15] NET050 NET049 NET037[0] 
+ NET037[1] NET037[2] NET037[3] NET037[4] NET037[5] NET037[6] NET037[7] 
+ NET037[8] NET037[9] NET037[10] NET037[11] NET037[12] NET037[13] NET037[14] 
+ NET037[15] NET039[0] NET039[1] NET039[2] NET039[3] NET039[4] NET039[5] 
+ NET039[6] NET039[7] NET039[8] NET039[9] NET039[10] NET039[11] NET039[12] 
+ NET039[13] NET039[14] NET039[15] NET052 NET051 NET048 NET047 NET045 NET046 
+ NET053 NET054 NET055 NET041 NET044[0] NET044[1] NET043[0] NET043[1] 
+ NET043[2] NET043[3] NET043[4] NET043[5] NET043[6] NET043[7] NET042[0] 
+ NET042[1] NET042[2] NET042[3] NET042[4] NET042[5] NET042[6] NET042[7] 
+ S1AHSF400W40_LIO_M16
XLIO_M8 NET057[0] NET057[1] NET057[2] NET057[3] NET057[4] NET057[5] NET057[6] 
+ NET057[7] NET056[0] NET056[1] NET056[2] NET056[3] NET056[4] NET056[5] 
+ NET056[6] NET056[7] NET069 NET068 NET059[0] NET059[1] NET059[2] NET059[3] 
+ NET059[4] NET059[5] NET059[6] NET059[7] NET058[0] NET058[1] NET058[2] 
+ NET058[3] NET058[4] NET058[5] NET058[6] NET058[7] NET071 NET070 NET067 
+ NET066 NET064 NET065 NET072 NET073 NET074 NET060 NET063[0] NET063[1] 
+ NET062[0] NET062[1] NET062[2] NET062[3] NET062[4] NET062[5] NET062[6] 
+ NET062[7] NET061[0] NET061[1] NET061[2] NET061[3] NET061[4] NET061[5] 
+ NET061[6] NET061[7] S1AHSF400W40_LIO_M8
XLIO_M4 NET50[0] NET50[1] NET50[2] NET50[3] NET49[0] NET49[1] NET49[2] 
+ NET49[3] NET46 NET45 NET52[0] NET52[1] NET52[2] NET52[3] NET51[0] NET51[1] 
+ NET51[2] NET51[3] NET48 NET47 NET44 NET43 NET41 NET42 NET53 NET54 NET55 
+ NET37 NET40[0] NET40[1] NET39[0] NET39[1] NET39[2] NET39[3] NET39[4] 
+ NET39[5] NET39[6] NET39[7] NET38[0] NET38[1] NET38[2] NET38[3] NET38[4] 
+ NET38[5] NET38[6] NET38[7] S1AHSF400W40_LIO_M4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    ARR_LIO_LD_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ARR_LIO_LD_SIM BLEQ_DN_LT BLEQ_DN_RT BLEQ_UP_LT BLEQ_UP_RT CVDDI RE_LT 
+ RE_RT SAEB_LT SAEB_RT VDDHD VDDI VSSI WE_LT WE_RT YL_LIO_LT[0] YL_LIO_LT[1] 
+ YL_LIO_RT[0] YL_LIO_RT[1] Y_DN_LT[0] Y_DN_LT[1] Y_DN_LT[2] Y_DN_LT[3] 
+ Y_DN_LT[4] Y_DN_LT[5] Y_DN_LT[6] Y_DN_LT[7] Y_DN_RT[0] Y_DN_RT[1] Y_DN_RT[2] 
+ Y_DN_RT[3] Y_DN_RT[4] Y_DN_RT[5] Y_DN_RT[6] Y_DN_RT[7] Y_UP_LT[0] Y_UP_LT[1] 
+ Y_UP_LT[2] Y_UP_LT[3] Y_UP_LT[4] Y_UP_LT[5] Y_UP_LT[6] Y_UP_LT[7] Y_UP_RT[0] 
+ Y_UP_RT[1] Y_UP_RT[2] Y_UP_RT[3] Y_UP_RT[4] Y_UP_RT[5] Y_UP_RT[6] Y_UP_RT[7]
*.PININFO BLEQ_DN_LT:B BLEQ_DN_RT:B BLEQ_UP_LT:B BLEQ_UP_RT:B CVDDI:B RE_LT:B 
*.PININFO RE_RT:B SAEB_LT:B SAEB_RT:B VDDHD:B VDDI:B VSSI:B WE_LT:B WE_RT:B 
*.PININFO YL_LIO_LT[0]:B YL_LIO_LT[1]:B YL_LIO_RT[0]:B YL_LIO_RT[1]:B 
*.PININFO Y_DN_LT[0]:B Y_DN_LT[1]:B Y_DN_LT[2]:B Y_DN_LT[3]:B Y_DN_LT[4]:B 
*.PININFO Y_DN_LT[5]:B Y_DN_LT[6]:B Y_DN_LT[7]:B Y_DN_RT[0]:B Y_DN_RT[1]:B 
*.PININFO Y_DN_RT[2]:B Y_DN_RT[3]:B Y_DN_RT[4]:B Y_DN_RT[5]:B Y_DN_RT[6]:B 
*.PININFO Y_DN_RT[7]:B Y_UP_LT[0]:B Y_UP_LT[1]:B Y_UP_LT[2]:B Y_UP_LT[3]:B 
*.PININFO Y_UP_LT[4]:B Y_UP_LT[5]:B Y_UP_LT[6]:B Y_UP_LT[7]:B Y_UP_RT[0]:B 
*.PININFO Y_UP_RT[1]:B Y_UP_RT[2]:B Y_UP_RT[3]:B Y_UP_RT[4]:B Y_UP_RT[5]:B 
*.PININFO Y_UP_RT[6]:B Y_UP_RT[7]:B
XLIO_M16 NET024[0] NET024[1] NET024[2] NET024[3] NET024[4] NET024[5] NET024[6] 
+ NET024[7] NET024[8] NET024[9] NET024[10] NET024[11] NET024[12] NET024[13] 
+ NET024[14] NET024[15] NET022[0] NET022[1] NET022[2] NET022[3] NET022[4] 
+ NET022[5] NET022[6] NET022[7] NET022[8] NET022[9] NET022[10] NET022[11] 
+ NET022[12] NET022[13] NET022[14] NET022[15] NET034 NET033 NET021[0] 
+ NET021[1] NET021[2] NET021[3] NET021[4] NET021[5] NET021[6] NET021[7] 
+ NET021[8] NET021[9] NET021[10] NET021[11] NET021[12] NET021[13] NET021[14] 
+ NET021[15] NET023[0] NET023[1] NET023[2] NET023[3] NET023[4] NET023[5] 
+ NET023[6] NET023[7] NET023[8] NET023[9] NET023[10] NET023[11] NET023[12] 
+ NET023[13] NET023[14] NET023[15] NET036 NET035 NET032 NET031 NET029 NET030 
+ NET037 NET038 NET039 NET025 NET028[0] NET028[1] NET027[0] NET027[1] 
+ NET027[2] NET027[3] NET027[4] NET027[5] NET027[6] NET027[7] NET026[0] 
+ NET026[1] NET026[2] NET026[3] NET026[4] NET026[5] NET026[6] NET026[7] 
+ S1AHSF400W40_LIO_M16
XLIO_M8 NET041[0] NET041[1] NET041[2] NET041[3] NET041[4] NET041[5] NET041[6] 
+ NET041[7] NET040[0] NET040[1] NET040[2] NET040[3] NET040[4] NET040[5] 
+ NET040[6] NET040[7] NET053 NET052 NET043[0] NET043[1] NET043[2] NET043[3] 
+ NET043[4] NET043[5] NET043[6] NET043[7] NET042[0] NET042[1] NET042[2] 
+ NET042[3] NET042[4] NET042[5] NET042[6] NET042[7] NET055 NET054 NET051 
+ NET050 NET048 NET049 NET056 NET057 NET058 NET044 NET047[0] NET047[1] 
+ NET046[0] NET046[1] NET046[2] NET046[3] NET046[4] NET046[5] NET046[6] 
+ NET046[7] NET045[0] NET045[1] NET045[2] NET045[3] NET045[4] NET045[5] 
+ NET045[6] NET045[7] S1AHSF400W40_LIO_M8
XLIO_M4 NET34[0] NET34[1] NET34[2] NET34[3] NET33[0] NET33[1] NET33[2] 
+ NET33[3] NET30 NET29 NET36[0] NET36[1] NET36[2] NET36[3] NET35[0] NET35[1] 
+ NET35[2] NET35[3] NET32 NET31 NET28 NET27 NET25 NET26 NET37 NET38 NET39 
+ NET21 NET24[0] NET24[1] NET23[0] NET23[1] NET23[2] NET23[3] NET23[4] 
+ NET23[5] NET23[6] NET23[7] NET22[0] NET22[1] NET22[2] NET22[3] NET22[4] 
+ NET22[5] NET22[6] NET22[7] S1AHSF400W40_LIO_M4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    TOP_EDGE
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TOP_EDGE VDDHD VDDI VSSI WLP_SAE WLP_SAE_TK
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B
XI248 WLP_SAE VSSI VDDHD NET54 S1AHSF400W40_AINV FN=1 WN=1.5U LN=0.06U FP=1 WP=2.5U 
+ LP=0.06U M=1
MM7 WLP_SAE_TK NET54 VSSI VSSI NCH L=60N W=3U M=2
MM3 WLP_SAE_TK NET54 VDDHD VDDI PCH L=60N W=4U M=2
MM0 WLP_SAE_TK NET54 VDDHD VDDI PCH L=60N W=2U M=2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_TOP_EDGE_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_TOP_EDGE_SIM VDDHD VDDI VSSI WLP_SAE_BT WLP_SAE_TK_BT
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE_BT:B WLP_SAE_TK_BT:B
XI1 NET09 NET08 NET010 NET06 NET07 S1AHSF400W40_TOP_EDGE
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    XDRV_LA512
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_XDRV_LA512 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] 
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] 
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WLOUT[0] WLOUT[1] WLPY 
+ WLPYB WLP_SAE WLP_SAE_TK YL[0]
*.PININFO DEC_Y[0]:I DEC_Y[1]:I DEC_Y[2]:I DEC_Y[3]:I DEC_Y[4]:I DEC_Y[5]:I 
*.PININFO DEC_Y[6]:I DEC_Y[7]:I PD_CVDDBUF:I WLPY:I WLPYB:I YL[0]:I WLOUT[0]:O 
*.PININFO WLOUT[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B PD_BUF:B RW_RE:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B
MM3 VDDI WLPY MWL2A VDDI PCH L=60N W=1U M=2
MP20 WLOUT[0] MWL2 VDDHD VDDI PCH L=60N W=4U M=4
MM5 MWL0A DEC_X1[0] VDDI VDDI PCH L=60N W=300N M=1
MM6 MWL0A DEC_X0[1] VDDI VDDI PCH L=60N W=300N M=1
MM0 MWL2A MWL1A VDDI VDDI PCH L=60N W=500N M=2
MM8 MWL2 MWL1 VDDI VDDI PCH L=60N W=500N M=2
MM1 WLOUT[1] MWL2A VDDHD VDDI PCH L=60N W=4U M=4
MP7 MWL0 DEC_X1[0] VDDI VDDI PCH L=60N W=300N M=1
MP4 VDDHD PD_BUF VDDI VDDI PCH L=60N W=2.5U M=4
MP6 MWL0 DEC_X0[0] VDDI VDDI PCH L=60N W=300N M=1
MP19 VDDI WLPY MWL2 VDDI PCH L=60N W=1U M=2
MP9 MWL0 DEC_X0[0] SH_NPD VSSI NCH L=60N W=300N M=1
MN6 WLOUT[0] MWL2 VSSI VSSI NCH L=60N W=4U M=2
MM7 MWL0A DEC_X0[1] SH_NPD VSSI NCH L=60N W=300N M=1
MN0 MWL2 MWL1 WLPYB VSSI NCH L=60N W=1.5U M=2
MM2 WLOUT[1] MWL2A VSSI VSSI NCH L=60N W=4U M=2
MM4 MWL2A MWL1A WLPYB VSSI NCH L=60N W=1.5U M=2
MN5 SH_NPD DEC_X1[0] VSSI VSSI NCH L=70N W=360.0N M=2
XINV1 MWL0 VSSI VDDHD MWL1 S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U LP=0.06U M=1
XI392 MWL0A VSSI VDDHD MWL1A S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U LP=0.06U 
+ M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    WLDV_2X1
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_WLDV_2X1 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[0] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI 
+ WL[0] WL[1] WL[2] WL[3] WLPY WLPYB WLP_SAE WLP_SAE_TK YL[0]
*.PININFO PD_BUF:I PD_CVDDBUF:I WLPY:I WLPYB:I DEC_X0[0]:B DEC_X0[1]:B 
*.PININFO DEC_X0[2]:B DEC_X0[3]:B DEC_X1[0]:B DEC_X2[0]:B DEC_X2[1]:B 
*.PININFO DEC_X2[2]:B DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B 
*.PININFO DEC_X3[3]:B DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B 
*.PININFO DEC_Y[0]:B DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B 
*.PININFO DEC_Y[6]:B DEC_Y[7]:B RW_RE:B VDDHD:B VDDI:B VSSI:B WL[0]:B WL[1]:B 
*.PININFO WL[2]:B WL[3]:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XWLDV_0 DEC_X0[0] DEC_X0[1] NET27[0] NET27[1] NET27[2] NET27[3] NET27[4] 
+ NET27[5] DEC_X1[0] NET25[0] NET25[1] NET25[2] NET25[3] NET25[4] NET25[5] 
+ NET25[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] 
+ DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] 
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD_BUF 
+ PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[0] WL[1] WLPY WLPYB WLP_SAE WLP_SAE_TK 
+ YL[0] S1AHSF400W40_XDRV_LA512
XWLDV_1 DEC_X0[2] DEC_X0[3] NET47[0] NET47[1] NET47[2] NET47[3] NET47[4] 
+ NET47[5] DEC_X1[0] NET45[0] NET45[1] NET45[2] NET45[3] NET45[4] NET45[5] 
+ NET45[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] 
+ DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] 
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] PD_BUF 
+ PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[2] WL[3] WLPY WLPYB WLP_SAE WLP_SAE_TK 
+ YL[0] S1AHSF400W40_XDRV_LA512
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_WLDV_LD_16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_WLDV_LD_16 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] 
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] PD_BUF VDDHD VDDI VSSI WLP_SAE WLP_SAE_TK YL[0]
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B DEC_X3[4]:B 
*.PININFO DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B DEC_Y[1]:B DEC_Y[2]:B 
*.PININFO DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B DEC_Y[7]:B PD_BUF:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XWLDV_2X1<2> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[1] NET035[0] 
+ NET035[1] NET035[2] NET035[3] NET034[0] NET034[1] NET034[2] NET034[3] 
+ NET034[4] NET034[5] NET034[6] NET034[7] NET033[0] NET033[1] NET033[2] 
+ NET033[3] NET033[4] NET033[5] NET033[6] NET033[7] PD_BUF NET021 NET032[0] 
+ VDDHD VDDI VSSI NET36[0] NET36[1] NET36[2] NET36[3] WLPY WLPYB NET031[0] 
+ NET030[0] NET029[0] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<3> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] NET035[4] 
+ NET035[5] NET035[6] NET035[7] NET034[8] NET034[9] NET034[10] NET034[11] 
+ NET034[12] NET034[13] NET034[14] NET034[15] NET033[8] NET033[9] NET033[10] 
+ NET033[11] NET033[12] NET033[13] NET033[14] NET033[15] PD_BUF NET021 
+ NET032[1] VDDHD VDDI VSSI NET36[4] NET36[5] NET36[6] NET36[7] WLPY WLPYB 
+ NET031[1] NET030[1] NET029[1] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<0> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[0] NET052[0] 
+ NET052[1] NET052[2] NET052[3] NET051[0] NET051[1] NET051[2] NET051[3] 
+ NET051[4] NET051[5] NET051[6] NET051[7] NET050[0] NET050[1] NET050[2] 
+ NET050[3] NET050[4] NET050[5] NET050[6] NET050[7] PD_BUF NET022 NET049[0] 
+ VDDHD VDDI VSSI NET46[0] NET46[1] NET46[2] NET46[3] WLPY WLPYB NET048[0] 
+ NET047[0] NET046[0] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<1> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] NET052[4] 
+ NET052[5] NET052[6] NET052[7] NET051[8] NET051[9] NET051[10] NET051[11] 
+ NET051[12] NET051[13] NET051[14] NET051[15] NET050[8] NET050[9] NET050[10] 
+ NET050[11] NET050[12] NET050[13] NET050[14] NET050[15] PD_BUF NET022 
+ NET049[1] VDDHD VDDI VSSI NET46[4] NET46[5] NET46[6] NET46[7] WLPY WLPYB 
+ NET048[1] NET047[1] NET046[1] S1AHSF400W40_WLDV_2X1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_WLDV_LD_32
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_WLDV_LD_32 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] 
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] PD_BUF VDDHD VDDI VSSI WLP_SAE WLP_SAE_TK YL[0]
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B DEC_X3[4]:B 
*.PININFO DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B DEC_Y[1]:B DEC_Y[2]:B 
*.PININFO DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B DEC_Y[7]:B PD_BUF:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XWLDV_2X1<2> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[1] NET040[0] 
+ NET040[1] NET040[2] NET040[3] NET039[0] NET039[1] NET039[2] NET039[3] 
+ NET039[4] NET039[5] NET039[6] NET039[7] NET038[0] NET038[1] NET038[2] 
+ NET038[3] NET038[4] NET038[5] NET038[6] NET038[7] PD_BUF NET021 NET037[0] 
+ VDDHD VDDI VSSI NET36[0] NET36[1] NET36[2] NET36[3] WLPY WLPYB NET036[0] 
+ NET035[0] NET034[0] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<3> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] NET040[4] 
+ NET040[5] NET040[6] NET040[7] NET039[8] NET039[9] NET039[10] NET039[11] 
+ NET039[12] NET039[13] NET039[14] NET039[15] NET038[8] NET038[9] NET038[10] 
+ NET038[11] NET038[12] NET038[13] NET038[14] NET038[15] PD_BUF NET021 
+ NET037[1] VDDHD VDDI VSSI NET36[4] NET36[5] NET36[6] NET36[7] WLPY WLPYB 
+ NET036[1] NET035[1] NET034[1] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<0> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[0] NET057[0] 
+ NET057[1] NET057[2] NET057[3] NET056[0] NET056[1] NET056[2] NET056[3] 
+ NET056[4] NET056[5] NET056[6] NET056[7] NET055[0] NET055[1] NET055[2] 
+ NET055[3] NET055[4] NET055[5] NET055[6] NET055[7] PD_BUF NET022 NET054[0] 
+ VDDHD VDDI VSSI NET46[0] NET46[1] NET46[2] NET46[3] WLPY WLPYB NET053[0] 
+ NET052[0] NET051[0] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<1> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] NET057[4] 
+ NET057[5] NET057[6] NET057[7] NET056[8] NET056[9] NET056[10] NET056[11] 
+ NET056[12] NET056[13] NET056[14] NET056[15] NET055[8] NET055[9] NET055[10] 
+ NET055[11] NET055[12] NET055[13] NET055[14] NET055[15] PD_BUF NET022 
+ NET054[1] VDDHD VDDI VSSI NET46[4] NET46[5] NET46[6] NET46[7] WLPY WLPYB 
+ NET053[1] NET052[1] NET051[1] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<6> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[3] NET074[0] 
+ NET074[1] NET074[2] NET074[3] NET073[0] NET073[1] NET073[2] NET073[3] 
+ NET073[4] NET073[5] NET073[6] NET073[7] NET072[0] NET072[1] NET072[2] 
+ NET072[3] NET072[4] NET072[5] NET072[6] NET072[7] PD_BUF NET016 NET071[0] 
+ VDDHD VDDI VSSI NET26[0] NET26[1] NET26[2] NET26[3] WLPY WLPYB NET070[0] 
+ NET069[0] NET068[0] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<7> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] NET074[4] 
+ NET074[5] NET074[6] NET074[7] NET073[8] NET073[9] NET073[10] NET073[11] 
+ NET073[12] NET073[13] NET073[14] NET073[15] NET072[8] NET072[9] NET072[10] 
+ NET072[11] NET072[12] NET072[13] NET072[14] NET072[15] PD_BUF NET016 
+ NET071[1] VDDHD VDDI VSSI NET26[4] NET26[5] NET26[6] NET26[7] WLPY WLPYB 
+ NET070[1] NET069[1] NET068[1] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<4> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[2] NET091[0] 
+ NET091[1] NET091[2] NET091[3] NET090[0] NET090[1] NET090[2] NET090[3] 
+ NET090[4] NET090[5] NET090[6] NET090[7] NET089[0] NET089[1] NET089[2] 
+ NET089[3] NET089[4] NET089[5] NET089[6] NET089[7] PD_BUF NET015 NET088[0] 
+ VDDHD VDDI VSSI NET16[0] NET16[1] NET16[2] NET16[3] WLPY WLPYB NET087[0] 
+ NET086[0] NET085[0] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<5> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] NET091[4] 
+ NET091[5] NET091[6] NET091[7] NET090[8] NET090[9] NET090[10] NET090[11] 
+ NET090[12] NET090[13] NET090[14] NET090[15] NET089[8] NET089[9] NET089[10] 
+ NET089[11] NET089[12] NET089[13] NET089[14] NET089[15] PD_BUF NET015 
+ NET088[1] VDDHD VDDI VSSI NET16[4] NET16[5] NET16[6] NET16[7] WLPY WLPYB 
+ NET087[1] NET086[1] NET085[1] S1AHSF400W40_WLDV_2X1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    WLDV_64X1
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_WLDV_64X1 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] PD_BUF PD_CVDDBUF VDDHD VDDI VSSI WL[0] WL[1] 
+ WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] 
+ WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] 
+ WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] 
+ WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] 
+ WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] 
+ WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] WLPY[0] WLPYB[0]
*.PININFO DEC_X0[0]:I DEC_X0[1]:I DEC_X0[2]:I DEC_X0[3]:I DEC_X0[4]:I 
*.PININFO DEC_X0[5]:I DEC_X0[6]:I DEC_X0[7]:I DEC_X1[0]:I DEC_X1[1]:I 
*.PININFO DEC_X1[2]:I DEC_X1[3]:I DEC_X1[4]:I DEC_X1[5]:I DEC_X1[6]:I 
*.PININFO DEC_X1[7]:I PD_BUF:I PD_CVDDBUF:I WLPY[0]:I WLPYB[0]:I WL[0]:O 
*.PININFO WL[1]:O WL[2]:O WL[3]:O WL[4]:O WL[5]:O WL[6]:O WL[7]:O WL[8]:O 
*.PININFO WL[9]:O WL[10]:O WL[11]:O WL[12]:O WL[13]:O WL[14]:O WL[15]:O 
*.PININFO WL[16]:O WL[17]:O WL[18]:O WL[19]:O WL[20]:O WL[21]:O WL[22]:O 
*.PININFO WL[23]:O WL[24]:O WL[25]:O WL[26]:O WL[27]:O WL[28]:O WL[29]:O 
*.PININFO WL[30]:O WL[31]:O WL[32]:O WL[33]:O WL[34]:O WL[35]:O WL[36]:O 
*.PININFO WL[37]:O WL[38]:O WL[39]:O WL[40]:O WL[41]:O WL[42]:O WL[43]:O 
*.PININFO WL[44]:O WL[45]:O WL[46]:O WL[47]:O WL[48]:O WL[49]:O WL[50]:O 
*.PININFO WL[51]:O WL[52]:O WL[53]:O WL[54]:O WL[55]:O WL[56]:O WL[57]:O 
*.PININFO WL[58]:O WL[59]:O WL[60]:O WL[61]:O WL[62]:O WL[63]:O VDDHD:B VDDI:B 
*.PININFO VSSI:B
XWLDV_2X1<0> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[0] NET17[0] 
+ NET17[1] NET17[2] NET17[3] NET16[0] NET16[1] NET16[2] NET16[3] NET16[4] 
+ NET16[5] NET16[6] NET16[7] NET15[0] NET15[1] NET15[2] NET15[3] NET15[4] 
+ NET15[5] NET15[6] NET15[7] PD_BUF PD_CVDDBUF NET14[0] VDDHD VDDI VSSI WL[0] 
+ WL[1] WL[2] WL[3] WLPY[0] WLPYB[0] NET13[0] NET12[0] NET11[0] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<1> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] NET17[4] 
+ NET17[5] NET17[6] NET17[7] NET16[8] NET16[9] NET16[10] NET16[11] NET16[12] 
+ NET16[13] NET16[14] NET16[15] NET15[8] NET15[9] NET15[10] NET15[11] 
+ NET15[12] NET15[13] NET15[14] NET15[15] PD_BUF PD_CVDDBUF NET14[1] VDDHD 
+ VDDI VSSI WL[4] WL[5] WL[6] WL[7] WLPY[0] WLPYB[0] NET13[1] NET12[1] 
+ NET11[1] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<2> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[1] NET17[8] 
+ NET17[9] NET17[10] NET17[11] NET16[16] NET16[17] NET16[18] NET16[19] 
+ NET16[20] NET16[21] NET16[22] NET16[23] NET15[16] NET15[17] NET15[18] 
+ NET15[19] NET15[20] NET15[21] NET15[22] NET15[23] PD_BUF PD_CVDDBUF NET14[2] 
+ VDDHD VDDI VSSI WL[8] WL[9] WL[10] WL[11] WLPY[0] WLPYB[0] NET13[2] NET12[2] 
+ NET11[2] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<3> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] NET17[12] 
+ NET17[13] NET17[14] NET17[15] NET16[24] NET16[25] NET16[26] NET16[27] 
+ NET16[28] NET16[29] NET16[30] NET16[31] NET15[24] NET15[25] NET15[26] 
+ NET15[27] NET15[28] NET15[29] NET15[30] NET15[31] PD_BUF PD_CVDDBUF NET14[3] 
+ VDDHD VDDI VSSI WL[12] WL[13] WL[14] WL[15] WLPY[0] WLPYB[0] NET13[3] 
+ NET12[3] NET11[3] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<4> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[2] NET17[16] 
+ NET17[17] NET17[18] NET17[19] NET16[32] NET16[33] NET16[34] NET16[35] 
+ NET16[36] NET16[37] NET16[38] NET16[39] NET15[32] NET15[33] NET15[34] 
+ NET15[35] NET15[36] NET15[37] NET15[38] NET15[39] PD_BUF PD_CVDDBUF NET14[4] 
+ VDDHD VDDI VSSI WL[16] WL[17] WL[18] WL[19] WLPY[0] WLPYB[0] NET13[4] 
+ NET12[4] NET11[4] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<5> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] NET17[20] 
+ NET17[21] NET17[22] NET17[23] NET16[40] NET16[41] NET16[42] NET16[43] 
+ NET16[44] NET16[45] NET16[46] NET16[47] NET15[40] NET15[41] NET15[42] 
+ NET15[43] NET15[44] NET15[45] NET15[46] NET15[47] PD_BUF PD_CVDDBUF NET14[5] 
+ VDDHD VDDI VSSI WL[20] WL[21] WL[22] WL[23] WLPY[0] WLPYB[0] NET13[5] 
+ NET12[5] NET11[5] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<6> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[3] NET17[24] 
+ NET17[25] NET17[26] NET17[27] NET16[48] NET16[49] NET16[50] NET16[51] 
+ NET16[52] NET16[53] NET16[54] NET16[55] NET15[48] NET15[49] NET15[50] 
+ NET15[51] NET15[52] NET15[53] NET15[54] NET15[55] PD_BUF PD_CVDDBUF NET14[6] 
+ VDDHD VDDI VSSI WL[24] WL[25] WL[26] WL[27] WLPY[0] WLPYB[0] NET13[6] 
+ NET12[6] NET11[6] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<7> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] NET17[28] 
+ NET17[29] NET17[30] NET17[31] NET16[56] NET16[57] NET16[58] NET16[59] 
+ NET16[60] NET16[61] NET16[62] NET16[63] NET15[56] NET15[57] NET15[58] 
+ NET15[59] NET15[60] NET15[61] NET15[62] NET15[63] PD_BUF PD_CVDDBUF NET14[7] 
+ VDDHD VDDI VSSI WL[28] WL[29] WL[30] WL[31] WLPY[0] WLPYB[0] NET13[7] 
+ NET12[7] NET11[7] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<8> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[4] NET17[32] 
+ NET17[33] NET17[34] NET17[35] NET16[64] NET16[65] NET16[66] NET16[67] 
+ NET16[68] NET16[69] NET16[70] NET16[71] NET15[64] NET15[65] NET15[66] 
+ NET15[67] NET15[68] NET15[69] NET15[70] NET15[71] PD_BUF PD_CVDDBUF NET14[8] 
+ VDDHD VDDI VSSI WL[32] WL[33] WL[34] WL[35] WLPY[0] WLPYB[0] NET13[8] 
+ NET12[8] NET11[8] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<9> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] NET17[36] 
+ NET17[37] NET17[38] NET17[39] NET16[72] NET16[73] NET16[74] NET16[75] 
+ NET16[76] NET16[77] NET16[78] NET16[79] NET15[72] NET15[73] NET15[74] 
+ NET15[75] NET15[76] NET15[77] NET15[78] NET15[79] PD_BUF PD_CVDDBUF NET14[9] 
+ VDDHD VDDI VSSI WL[36] WL[37] WL[38] WL[39] WLPY[0] WLPYB[0] NET13[9] 
+ NET12[9] NET11[9] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<10> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[5] NET17[40] 
+ NET17[41] NET17[42] NET17[43] NET16[80] NET16[81] NET16[82] NET16[83] 
+ NET16[84] NET16[85] NET16[86] NET16[87] NET15[80] NET15[81] NET15[82] 
+ NET15[83] NET15[84] NET15[85] NET15[86] NET15[87] PD_BUF PD_CVDDBUF 
+ NET14[10] VDDHD VDDI VSSI WL[40] WL[41] WL[42] WL[43] WLPY[0] WLPYB[0] 
+ NET13[10] NET12[10] NET11[10] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<11> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] NET17[44] 
+ NET17[45] NET17[46] NET17[47] NET16[88] NET16[89] NET16[90] NET16[91] 
+ NET16[92] NET16[93] NET16[94] NET16[95] NET15[88] NET15[89] NET15[90] 
+ NET15[91] NET15[92] NET15[93] NET15[94] NET15[95] PD_BUF PD_CVDDBUF 
+ NET14[11] VDDHD VDDI VSSI WL[44] WL[45] WL[46] WL[47] WLPY[0] WLPYB[0] 
+ NET13[11] NET12[11] NET11[11] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<12> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[6] NET17[48] 
+ NET17[49] NET17[50] NET17[51] NET16[96] NET16[97] NET16[98] NET16[99] 
+ NET16[100] NET16[101] NET16[102] NET16[103] NET15[96] NET15[97] NET15[98] 
+ NET15[99] NET15[100] NET15[101] NET15[102] NET15[103] PD_BUF PD_CVDDBUF 
+ NET14[12] VDDHD VDDI VSSI WL[48] WL[49] WL[50] WL[51] WLPY[0] WLPYB[0] 
+ NET13[12] NET12[12] NET11[12] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<13> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] NET17[52] 
+ NET17[53] NET17[54] NET17[55] NET16[104] NET16[105] NET16[106] NET16[107] 
+ NET16[108] NET16[109] NET16[110] NET16[111] NET15[104] NET15[105] NET15[106] 
+ NET15[107] NET15[108] NET15[109] NET15[110] NET15[111] PD_BUF PD_CVDDBUF 
+ NET14[13] VDDHD VDDI VSSI WL[52] WL[53] WL[54] WL[55] WLPY[0] WLPYB[0] 
+ NET13[13] NET12[13] NET11[13] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<14> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[7] NET17[56] 
+ NET17[57] NET17[58] NET17[59] NET16[112] NET16[113] NET16[114] NET16[115] 
+ NET16[116] NET16[117] NET16[118] NET16[119] NET15[112] NET15[113] NET15[114] 
+ NET15[115] NET15[116] NET15[117] NET15[118] NET15[119] PD_BUF PD_CVDDBUF 
+ NET14[14] VDDHD VDDI VSSI WL[56] WL[57] WL[58] WL[59] WLPY[0] WLPYB[0] 
+ NET13[14] NET12[14] NET11[14] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<15> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] NET17[60] 
+ NET17[61] NET17[62] NET17[63] NET16[120] NET16[121] NET16[122] NET16[123] 
+ NET16[124] NET16[125] NET16[126] NET16[127] NET15[120] NET15[121] NET15[122] 
+ NET15[123] NET15[124] NET15[125] NET15[126] NET15[127] PD_BUF PD_CVDDBUF 
+ NET14[15] VDDHD VDDI VSSI WL[60] WL[61] WL[62] WL[63] WLPY[0] WLPYB[0] 
+ NET13[15] NET12[15] NET11[15] S1AHSF400W40_WLDV_2X1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_WLDV_LD_64
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_WLDV_LD_64 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] 
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] PD_BUF VDDHD VDDI VSSI WLP_SAE WLP_SAE_TK YL[0]
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B DEC_X3[4]:B 
*.PININFO DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B DEC_Y[1]:B DEC_Y[2]:B 
*.PININFO DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B DEC_Y[7]:B PD_BUF:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XI28 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] PD_BUF NET34 VDDHD VDDI VSSI NET30[0] NET30[1] NET30[2] 
+ NET30[3] NET30[4] NET30[5] NET30[6] NET30[7] NET30[8] NET30[9] NET30[10] 
+ NET30[11] NET30[12] NET30[13] NET30[14] NET30[15] NET30[16] NET30[17] 
+ NET30[18] NET30[19] NET30[20] NET30[21] NET30[22] NET30[23] NET30[24] 
+ NET30[25] NET30[26] NET30[27] NET30[28] NET30[29] NET30[30] NET30[31] 
+ NET30[32] NET30[33] NET30[34] NET30[35] NET30[36] NET30[37] NET30[38] 
+ NET30[39] NET30[40] NET30[41] NET30[42] NET30[43] NET30[44] NET30[45] 
+ NET30[46] NET30[47] NET30[48] NET30[49] NET30[50] NET30[51] NET30[52] 
+ NET30[53] NET30[54] NET30[55] NET30[56] NET30[57] NET30[58] NET30[59] 
+ NET30[60] NET30[61] NET30[62] NET30[63] NET26 NET25 S1AHSF400W40_WLDV_64X1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    XDRV_STRAP
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_XDRV_STRAP VDDHD VDDI VSSI WLPY WLPYB
*.PININFO WLPY:I VDDHD:B VDDI:B VSSI:B WLPYB:B
MP0 WLPYB WLPY VDDHD VDDI PCH L=60N W=3U M=2
MN1 WLPYB WLPY VSSI VSSI NCH L=60N W=4U M=2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_WLDV_LD_128
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_WLDV_LD_128 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] 
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] PD_BUF VDDHD VDDI VSSI WLP_SAE WLP_SAE_TK YL[0]
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B DEC_X3[4]:B 
*.PININFO DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B DEC_Y[1]:B DEC_Y[2]:B 
*.PININFO DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B DEC_Y[7]:B PD_BUF:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XI28 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] PD_BUF NET071 VDDHD VDDI VSSI NET35[0] NET35[1] NET35[2] 
+ NET35[3] NET35[4] NET35[5] NET35[6] NET35[7] NET35[8] NET35[9] NET35[10] 
+ NET35[11] NET35[12] NET35[13] NET35[14] NET35[15] NET35[16] NET35[17] 
+ NET35[18] NET35[19] NET35[20] NET35[21] NET35[22] NET35[23] NET35[24] 
+ NET35[25] NET35[26] NET35[27] NET35[28] NET35[29] NET35[30] NET35[31] 
+ NET35[32] NET35[33] NET35[34] NET35[35] NET35[36] NET35[37] NET35[38] 
+ NET35[39] NET35[40] NET35[41] NET35[42] NET35[43] NET35[44] NET35[45] 
+ NET35[46] NET35[47] NET35[48] NET35[49] NET35[50] NET35[51] NET35[52] 
+ NET35[53] NET35[54] NET35[55] NET35[56] NET35[57] NET35[58] NET35[59] 
+ NET35[60] NET35[61] NET35[62] NET35[63] NET31 NET30 S1AHSF400W40_WLDV_64X1
XI25 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] PD_BUF NET061 VDDHD VDDI VSSI NET45[0] NET45[1] NET45[2] 
+ NET45[3] NET45[4] NET45[5] NET45[6] NET45[7] NET45[8] NET45[9] NET45[10] 
+ NET45[11] NET45[12] NET45[13] NET45[14] NET45[15] NET45[16] NET45[17] 
+ NET45[18] NET45[19] NET45[20] NET45[21] NET45[22] NET45[23] NET45[24] 
+ NET45[25] NET45[26] NET45[27] NET45[28] NET45[29] NET45[30] NET45[31] 
+ NET45[32] NET45[33] NET45[34] NET45[35] NET45[36] NET45[37] NET45[38] 
+ NET45[39] NET45[40] NET45[41] NET45[42] NET45[43] NET45[44] NET45[45] 
+ NET45[46] NET45[47] NET45[48] NET45[49] NET45[50] NET45[51] NET45[52] 
+ NET45[53] NET45[54] NET45[55] NET45[56] NET45[57] NET45[58] NET45[59] 
+ NET45[60] NET45[61] NET45[62] NET45[63] NET039 NET038 S1AHSF400W40_WLDV_64X1
XI24 VDDHD VDDI VSSI NET063 NET065 S1AHSF400W40_XDRV_STRAP
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_WLDV_LD_256
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_WLDV_LD_256 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] 
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] PD_BUF VDDHD VDDI VSSI WLP_SAE WLP_SAE_TK YL[0]
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B DEC_X3[4]:B 
*.PININFO DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B DEC_Y[1]:B DEC_Y[2]:B 
*.PININFO DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B DEC_Y[7]:B PD_BUF:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XI28 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] PD_BUF NET071 VDDHD VDDI VSSI NET35[0] NET35[1] NET35[2] 
+ NET35[3] NET35[4] NET35[5] NET35[6] NET35[7] NET35[8] NET35[9] NET35[10] 
+ NET35[11] NET35[12] NET35[13] NET35[14] NET35[15] NET35[16] NET35[17] 
+ NET35[18] NET35[19] NET35[20] NET35[21] NET35[22] NET35[23] NET35[24] 
+ NET35[25] NET35[26] NET35[27] NET35[28] NET35[29] NET35[30] NET35[31] 
+ NET35[32] NET35[33] NET35[34] NET35[35] NET35[36] NET35[37] NET35[38] 
+ NET35[39] NET35[40] NET35[41] NET35[42] NET35[43] NET35[44] NET35[45] 
+ NET35[46] NET35[47] NET35[48] NET35[49] NET35[50] NET35[51] NET35[52] 
+ NET35[53] NET35[54] NET35[55] NET35[56] NET35[57] NET35[58] NET35[59] 
+ NET35[60] NET35[61] NET35[62] NET35[63] NET31 NET30 S1AHSF400W40_WLDV_64X1
XWLDV_64X1_0 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] PD_BUF NET041 VDDHD VDDI VSSI NET19[0] 
+ NET19[1] NET19[2] NET19[3] NET19[4] NET19[5] NET19[6] NET19[7] NET19[8] 
+ NET19[9] NET19[10] NET19[11] NET19[12] NET19[13] NET19[14] NET19[15] 
+ NET19[16] NET19[17] NET19[18] NET19[19] NET19[20] NET19[21] NET19[22] 
+ NET19[23] NET19[24] NET19[25] NET19[26] NET19[27] NET19[28] NET19[29] 
+ NET19[30] NET19[31] NET19[32] NET19[33] NET19[34] NET19[35] NET19[36] 
+ NET19[37] NET19[38] NET19[39] NET19[40] NET19[41] NET19[42] NET19[43] 
+ NET19[44] NET19[45] NET19[46] NET19[47] NET19[48] NET19[49] NET19[50] 
+ NET19[51] NET19[52] NET19[53] NET19[54] NET19[55] NET19[56] NET19[57] 
+ NET19[58] NET19[59] NET19[60] NET19[61] NET19[62] NET19[63] NET029 NET028 
+ S1AHSF400W40_WLDV_64X1
XI25 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] PD_BUF NET061 VDDHD VDDI VSSI NET45[0] NET45[1] NET45[2] 
+ NET45[3] NET45[4] NET45[5] NET45[6] NET45[7] NET45[8] NET45[9] NET45[10] 
+ NET45[11] NET45[12] NET45[13] NET45[14] NET45[15] NET45[16] NET45[17] 
+ NET45[18] NET45[19] NET45[20] NET45[21] NET45[22] NET45[23] NET45[24] 
+ NET45[25] NET45[26] NET45[27] NET45[28] NET45[29] NET45[30] NET45[31] 
+ NET45[32] NET45[33] NET45[34] NET45[35] NET45[36] NET45[37] NET45[38] 
+ NET45[39] NET45[40] NET45[41] NET45[42] NET45[43] NET45[44] NET45[45] 
+ NET45[46] NET45[47] NET45[48] NET45[49] NET45[50] NET45[51] NET45[52] 
+ NET45[53] NET45[54] NET45[55] NET45[56] NET45[57] NET45[58] NET45[59] 
+ NET45[60] NET45[61] NET45[62] NET45[63] NET039 NET038 S1AHSF400W40_WLDV_64X1
XI27 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] PD_BUF NET051 VDDHD VDDI VSSI NET18[0] NET18[1] NET18[2] 
+ NET18[3] NET18[4] NET18[5] NET18[6] NET18[7] NET18[8] NET18[9] NET18[10] 
+ NET18[11] NET18[12] NET18[13] NET18[14] NET18[15] NET18[16] NET18[17] 
+ NET18[18] NET18[19] NET18[20] NET18[21] NET18[22] NET18[23] NET18[24] 
+ NET18[25] NET18[26] NET18[27] NET18[28] NET18[29] NET18[30] NET18[31] 
+ NET18[32] NET18[33] NET18[34] NET18[35] NET18[36] NET18[37] NET18[38] 
+ NET18[39] NET18[40] NET18[41] NET18[42] NET18[43] NET18[44] NET18[45] 
+ NET18[46] NET18[47] NET18[48] NET18[49] NET18[50] NET18[51] NET18[52] 
+ NET18[53] NET18[54] NET18[55] NET18[56] NET18[57] NET18[58] NET18[59] 
+ NET18[60] NET18[61] NET18[62] NET18[63] NET049 NET048 S1AHSF400W40_WLDV_64X1
XXDRV_STRP_0 VDDHD VDDI VSSI NET058 NET060 S1AHSF400W40_XDRV_STRAP
XI24 VDDHD VDDI VSSI NET063 NET065 S1AHSF400W40_XDRV_STRAP
XI26 VDDHD VDDI VSSI NET068 NET070 S1AHSF400W40_XDRV_STRAP
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_WLDV_LD_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_WLDV_LD_SIM CVDDHD CVDDI DEC_X0_BT[0] DEC_X0_BT[1] DEC_X0_BT[2] 
+ DEC_X0_BT[3] DEC_X0_BT[4] DEC_X0_BT[5] DEC_X0_BT[6] DEC_X0_BT[7] 
+ DEC_X0_TP[0] DEC_X0_TP[1] DEC_X0_TP[2] DEC_X0_TP[3] DEC_X0_TP[4] 
+ DEC_X0_TP[5] DEC_X0_TP[6] DEC_X0_TP[7] DEC_X1_BT[0] DEC_X1_BT[1] 
+ DEC_X1_BT[2] DEC_X1_BT[3] DEC_X1_BT[4] DEC_X1_BT[5] DEC_X1_BT[6] 
+ DEC_X1_BT[7] DEC_X1_TP[0] DEC_X1_TP[1] DEC_X1_TP[2] DEC_X1_TP[3] 
+ DEC_X1_TP[4] DEC_X1_TP[5] DEC_X1_TP[6] DEC_X1_TP[7] DEC_X2_BT[0] 
+ DEC_X2_BT[1] DEC_X2_BT[2] DEC_X2_BT[3] DEC_X2_TP[0] DEC_X2_TP[1] 
+ DEC_X2_TP[2] DEC_X2_TP[3] DEC_X3_BT[0] DEC_X3_BT[1] DEC_X3_BT[2] 
+ DEC_X3_BT[3] DEC_X3_BT[4] DEC_X3_BT[5] DEC_X3_BT[6] DEC_X3_BT[7] 
+ DEC_X3_TP[0] DEC_X3_TP[1] DEC_X3_TP[2] DEC_X3_TP[3] DEC_X3_TP[4] 
+ DEC_X3_TP[5] DEC_X3_TP[6] DEC_X3_TP[7] DEC_Y_BT[0] DEC_Y_BT[1] DEC_Y_BT[2] 
+ DEC_Y_BT[3] DEC_Y_BT[4] DEC_Y_BT[5] DEC_Y_BT[6] DEC_Y_BT[7] DEC_Y_TP[0] 
+ DEC_Y_TP[1] DEC_Y_TP[2] DEC_Y_TP[3] DEC_Y_TP[4] DEC_Y_TP[5] DEC_Y_TP[6] 
+ DEC_Y_TP[7] PD_BUF_BT PD_BUF_TP PD_CVDDBUF_BT PD_CVDDBUF_TP RW_RE_BT 
+ RW_RE_TP VDDHD VDDI VSSI WLP_SAE_BT WLP_SAE_TK_BT WLP_SAE_TK_TP WLP_SAE_TP 
+ YL_BT[0] YL_TP[0]
*.PININFO DEC_X0_BT[0]:I DEC_X0_BT[1]:I DEC_X0_BT[2]:I DEC_X0_BT[3]:I 
*.PININFO DEC_X0_BT[4]:I DEC_X0_BT[5]:I DEC_X0_BT[6]:I DEC_X0_BT[7]:I 
*.PININFO DEC_X1_BT[0]:I DEC_X1_BT[1]:I DEC_X1_BT[2]:I DEC_X1_BT[3]:I 
*.PININFO DEC_X1_BT[4]:I DEC_X1_BT[5]:I DEC_X1_BT[6]:I DEC_X1_BT[7]:I 
*.PININFO PD_BUF_BT:I PD_CVDDBUF_BT:I RW_RE_TP:I DEC_X0_TP[0]:O DEC_X0_TP[1]:O 
*.PININFO DEC_X0_TP[2]:O DEC_X0_TP[3]:O DEC_X0_TP[4]:O DEC_X0_TP[5]:O 
*.PININFO DEC_X0_TP[6]:O DEC_X0_TP[7]:O DEC_X1_TP[0]:O DEC_X1_TP[1]:O 
*.PININFO DEC_X1_TP[2]:O DEC_X1_TP[3]:O DEC_X1_TP[4]:O DEC_X1_TP[5]:O 
*.PININFO DEC_X1_TP[6]:O DEC_X1_TP[7]:O PD_BUF_TP:O PD_CVDDBUF_TP:O CVDDHD:B 
*.PININFO CVDDI:B DEC_X2_BT[0]:B DEC_X2_BT[1]:B DEC_X2_BT[2]:B DEC_X2_BT[3]:B 
*.PININFO DEC_X2_TP[0]:B DEC_X2_TP[1]:B DEC_X2_TP[2]:B DEC_X2_TP[3]:B 
*.PININFO DEC_X3_BT[0]:B DEC_X3_BT[1]:B DEC_X3_BT[2]:B DEC_X3_BT[3]:B 
*.PININFO DEC_X3_BT[4]:B DEC_X3_BT[5]:B DEC_X3_BT[6]:B DEC_X3_BT[7]:B 
*.PININFO DEC_X3_TP[0]:B DEC_X3_TP[1]:B DEC_X3_TP[2]:B DEC_X3_TP[3]:B 
*.PININFO DEC_X3_TP[4]:B DEC_X3_TP[5]:B DEC_X3_TP[6]:B DEC_X3_TP[7]:B 
*.PININFO DEC_Y_BT[0]:B DEC_Y_BT[1]:B DEC_Y_BT[2]:B DEC_Y_BT[3]:B 
*.PININFO DEC_Y_BT[4]:B DEC_Y_BT[5]:B DEC_Y_BT[6]:B DEC_Y_BT[7]:B 
*.PININFO DEC_Y_TP[0]:B DEC_Y_TP[1]:B DEC_Y_TP[2]:B DEC_Y_TP[3]:B 
*.PININFO DEC_Y_TP[4]:B DEC_Y_TP[5]:B DEC_Y_TP[6]:B DEC_Y_TP[7]:B RW_RE_BT:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE_BT:B WLP_SAE_TK_BT:B WLP_SAE_TK_TP:B 
*.PININFO WLP_SAE_TP:B YL_BT[0]:B YL_TP[0]:B
XI38 NET09[0] NET09[1] NET09[2] NET09[3] NET09[4] NET09[5] NET09[6] NET09[7] 
+ NET010[0] NET010[1] NET010[2] NET010[3] NET010[4] NET010[5] NET010[6] 
+ NET010[7] NET06[0] NET06[1] NET06[2] NET06[3] NET012[0] NET012[1] NET012[2] 
+ NET012[3] NET012[4] NET012[5] NET012[6] NET012[7] NET011[0] NET011[1] 
+ NET011[2] NET011[3] NET011[4] NET011[5] NET011[6] NET011[7] NET05 NET042 
+ NET041 NET043 NET07 NET040 NET08 S1AHSF400W40_BK_WLDV_LD_16
XI39 NET049[0] NET049[1] NET049[2] NET049[3] NET049[4] NET049[5] NET049[6] 
+ NET049[7] NET048[0] NET048[1] NET048[2] NET048[3] NET048[4] NET048[5] 
+ NET048[6] NET048[7] NET047[0] NET047[1] NET047[2] NET047[3] NET046[0] 
+ NET046[1] NET046[2] NET046[3] NET046[4] NET046[5] NET046[6] NET046[7] 
+ NET050[0] NET050[1] NET050[2] NET050[3] NET050[4] NET050[5] NET050[6] 
+ NET050[7] NET044 NET054 NET053 NET055 NET051 NET052 NET045 S1AHSF400W40_BK_WLDV_LD_32
XI34 NET40[0] NET40[1] NET40[2] NET40[3] NET40[4] NET40[5] NET40[6] NET40[7] 
+ NET36[0] NET36[1] NET36[2] NET36[3] NET36[4] NET36[5] NET36[6] NET36[7] 
+ NET35[0] NET35[1] NET35[2] NET35[3] NET34[0] NET34[1] NET34[2] NET34[3] 
+ NET34[4] NET34[5] NET34[6] NET34[7] NET031[0] NET031[1] NET031[2] NET031[3] 
+ NET031[4] NET031[5] NET031[6] NET031[7] NET32 NET42 NET41 NET43 NET030 
+ NET029 NET028 S1AHSF400W40_BK_WLDV_LD_64
XI35 NET033[0] NET033[1] NET033[2] NET033[3] NET033[4] NET033[5] NET033[6] 
+ NET033[7] NET032[0] NET032[1] NET032[2] NET032[3] NET032[4] NET032[5] 
+ NET032[6] NET032[7] NET01[0] NET01[1] NET01[2] NET01[3] NET04[0] NET04[1] 
+ NET04[2] NET04[3] NET04[4] NET04[5] NET04[6] NET04[7] NET034[0] NET034[1] 
+ NET034[2] NET034[3] NET034[4] NET034[5] NET034[6] NET034[7] NET03 NET038 
+ NET037 NET039 NET035 NET036 NET02 S1AHSF400W40_BK_WLDV_LD_128
XI36 NET085[0] NET085[1] NET085[2] NET085[3] NET085[4] NET085[5] NET085[6] 
+ NET085[7] NET084[0] NET084[1] NET084[2] NET084[3] NET084[4] NET084[5] 
+ NET084[6] NET084[7] NET083[0] NET083[1] NET083[2] NET083[3] NET082[0] 
+ NET082[1] NET082[2] NET082[3] NET082[4] NET082[5] NET082[6] NET082[7] 
+ NET086[0] NET086[1] NET086[2] NET086[3] NET086[4] NET086[5] NET086[6] 
+ NET086[7] NET080 NET090 NET089 NET091 NET087 NET088 NET081 S1AHSF400W40_BK_WLDV_LD_256
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    XDRV_WLP_F
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_XDRV_WLP_F BLEQ BLEQB BS PD_BUF RD_RST VDDHD VDDI VSSI WLOUT
*.PININFO BS:I PD_BUF:I RD_RST:I BLEQ:O BLEQB:O WLOUT:O VDDHD:B VDDI:B VSSI:B
XI235 BS NET102 VSSI VDDHD MWL S1AHSF400W40_ANAND FN2=2 WN2=1.5U LN2=0.06U FN1=2 WN1=1.5U 
+ LN1=0.06U FP1=2 WP1=1.5U LP1=0.06U FP2=2 WP2=1.5U LP2=0.06U M=1
XI530 BS D3 VSSI VDDHD NET78 S1AHSF400W40_ANAND FN2=2 WN2=1.5U LN2=0.06U FN1=2 WN1=1.5U 
+ LN1=0.06U FP1=2 WP1=1.5U LP1=0.06U FP2=2 WP2=1.5U LP2=0.06U M=1
MM0 BLEQB PD_BUF VSSI VSSI NCH L=60N W=1U M=1
XI527 MWL VSSI VDDHD WLOUT S1AHSF400W40_AINV FN=6 WN=1U LN=0.06U FP=6 WP=2U LP=0.06U M=1
XI507 RD_RST VSSI VDDHD D1 S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.6U LP=0.06U 
+ M=1
XI539 BLEQB VSSI VDDI BLEQ S1AHSF400W40_AINV FN=16 WN=1.5U LN=0.07U FP=16 WP=3U LP=0.07U 
+ M=1
XI522 D3 VSSI VDDHD D4 S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.6U LP=0.06U M=1
XI521 D2 VSSI VDDHD D3 S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.6U LP=0.06U M=1
XI520 D1 VSSI VDDHD D2 S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.6U LP=0.06U M=1
XI538 NET78 VSSI VDDHD BLEQB S1AHSF400W40_AINV FN=6 WN=1U LN=0.06U FP=6 WP=2U LP=0.06U M=1
XI529 RD_RST VSSI VDDHD NET102 S1AHSF400W40_AINV FN=1 WN=0.4U LN=0.06U FP=1 WP=0.8U 
+ LP=0.06U M=1
XI533 D4 VSSI VDDHD D5 S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.6U LP=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65_LOGIC
* CELL NAME:    NAND_BULK
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_NAND_BULK A B G GB P PB Y
*.PININFO A:I B:I G:I GB:I P:I PB:I Y:O
M1 Y B P PB PCH L=LP2 W=WP2 M=1*FP2
M4 Y A P PB PCH L=LP1 W=WP1 M=1*FP1
M6 NET9 A G GB NCH L=LN1 W=WN1 M=1*FN1
M8 Y B NET9 GB NCH L=LN2 W=WN2 M=1*FN2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    XDRV_READ
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_XDRV_READ BS PD_BUF SAEB VDDHD VDDI VSSI WLP_SAE
*.PININFO BS:I PD_BUF:I WLP_SAE:I SAEB:O VDDHD:B VDDI:B VSSI:B
XI424 BS WLP_SAE VSSI VSSI VDDHD VDDI BS_WLPSAEB S1AHSF400W40_NAND_BULK FN2=1 WN2=1.2U 
+ LN2=0.06U FN1=1 WN1=1.2U LN1=0.06U FP1=1 WP1=1.2U LP1=0.06U FP2=1 WP2=1.2U 
+ LP2=0.06U M=1
MP19 SAEB BS_WLPSAEB VDDHD VDDI PCH L=60N W=1.2U M=4
MN1 SAEB PD_BUF VSSI VSSI NCH L=60N W=600N M=1
MN20 SAEB BS_WLPSAEB VSSI VSSI NCH L=60N W=1.2U M=2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    XDRV_Y10
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_XDRV_Y10 BSB PD_BUF VDDHD VSSI YIN YOUT[0] YOUT[1]
*.PININFO BSB:I PD_BUF:I YIN:I YOUT[0]:O YOUT[1]:O VDDHD:B VSSI:B
XI381 BSB VSSI VDDHD BSB1B S1AHSF400W40_AINV FN=1 WN=0.8U LN=0.06U FP=1 WP=1.6U LP=0.06U 
+ M=1
XI25 YINL VSSI VDDHD YINL1B S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U LP=0.06U 
+ M=1
XI383 YINL1B BSB1B VSSI VDDHD NET112 S1AHSF400W40_ANAND FN2=1 WN2=1.5U LN2=0.06U FN1=1 
+ WN1=1.5U LN1=0.06U FP1=1 WP1=1.5U LP1=0.06U FP2=1 WP2=1.5U LP2=0.06U M=2
XNAND0 YINL BSB1B VSSI VDDHD NET107 S1AHSF400W40_ANAND FN2=1 WN2=1.5U LN2=0.06U FN1=1 
+ WN1=1.5U LN1=0.06U FP1=1 WP1=1.5U LP1=0.06U FP2=1 WP2=1.5U LP2=0.06U M=2
MM19 YINL YIN N7 VSSI NCH L=60N W=1U M=1
MM20 YINL BSB1B NET136 VSSI NCH L=60N W=300N M=1
MM21 NET136 YINL1B VSSI VSSI NCH L=60N W=300N M=1
MM23 N7 BSB VSSI VSSI NCH L=60N W=1U M=1
MM0 YOUT[0] PD_BUF VSSI VSSI NCH L=60N W=150.0N M=4
MM3 YOUT[1] PD_BUF VSSI VSSI NCH L=60N W=150.0N M=4
MN19 YOUT[0] NET107 VSSI VSSI NCH L=60N W=1.5U M=4
MM2 YOUT[1] NET112 VSSI VSSI NCH L=60N W=1.5U M=4
MM26 YINL BSB NET171 VDDHD PCH L=60N W=500N M=1
MP28 YOUT[0] NET107 VDDHD VDDHD PCH L=60N W=3U M=4
MM27 NET171 YINL1B VDDHD VDDHD PCH L=60N W=500N M=1
MM28 N5 BSB1B VDDHD VDDHD PCH L=60N W=1U M=2
MM29 YINL YIN N5 VDDHD PCH L=60N W=1U M=2
MM1 YOUT[1] NET112 VDDHD VDDHD PCH L=60N W=3U M=4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    XDRV_RW
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_XDRV_RW BS PD_BUF RE VDDHD VSSI WE WLP
*.PININFO BS:I PD_BUF:I WLP:I RE:O WE:O VDDHD:B VSSI:B
MN17 WE PD_BUF VSSI VSSI NCH L=60N W=150.0N M=4
MN3 RE PD_BUF VSSI VSSI NCH L=60N W=150.0N M=4
XINV0 Z0 VSSI VDDHD RE S1AHSF400W40_AINV FN=1 WN=1.5U LN=0.06U FP=1 WP=3U LP=0.06U M=4
XINV1 Z0 VSSI VDDHD Z1 S1AHSF400W40_AINV FN=1 WN=0.62U LN=0.06U FP=1 WP=1.25U LP=0.06U M=2
XINV2 Z1 VSSI VDDHD WE S1AHSF400W40_AINV FN=1 WN=1.5U LN=0.06U FP=1 WP=3U LP=0.06U M=4
XNAND0 WLP BS VSSI VDDHD Z0 S1AHSF400W40_ANAND FN2=2 WN2=1.25U LN2=0.06U FN1=2 WN1=1.25U 
+ LN1=0.06U FP1=2 WP1=1.25U LP1=0.06U FP2=2 WP2=1.25U LP2=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    XDRV_Y4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_XDRV_Y4 PD_BUF VDDHD VSSI WLPY YIN[0] YIN[1] YIN[2] YIN[3] YOUT[0] 
+ YOUT[1] YOUT[2] YOUT[3]
*.PININFO PD_BUF:I WLPY:I YIN[0]:I YIN[1]:I YIN[2]:I YIN[3]:I YOUT[0]:O 
*.PININFO YOUT[1]:O YOUT[2]:O YOUT[3]:O VDDHD:B VSSI:B
MM9 YOUT[2] MWL2[2] VDDHD VDDHD PCH L=60N W=3U M=4
MM10 MWL2[2] WLPY VDDHD VDDHD PCH L=60N W=750.0N M=4
MM12 MWL2[2] YIN[2] VDDHD VDDHD PCH L=60N W=750.0N M=4
MM13 MWL2[3] YIN[3] VDDHD VDDHD PCH L=60N W=750.0N M=4
MM15 MWL2[3] WLPY VDDHD VDDHD PCH L=60N W=750.0N M=4
MM16 YOUT[3] MWL2[3] VDDHD VDDHD PCH L=60N W=3U M=4
MM3 MWL2[1] YIN[1] VDDHD VDDHD PCH L=60N W=750.0N M=4
MP28 YOUT[0] MWL2[0] VDDHD VDDHD PCH L=60N W=3U M=4
MP31 SHARE WLPY VDDHD VDDHD PCH L=60N W=750.0N M=1
MP16 MWL2[0] YIN[0] VDDHD VDDHD PCH L=60N W=750.0N M=4
MM5 MWL2[1] WLPY VDDHD VDDHD PCH L=60N W=750.0N M=4
MM6 YOUT[1] MWL2[1] VDDHD VDDHD PCH L=60N W=3U M=4
MP30 MWL2[0] WLPY VDDHD VDDHD PCH L=60N W=750.0N M=4
MM11 MWL2[2] YIN[2] SHARE VSSI NCH L=60N W=1.5U M=4
MM14 MWL2[3] YIN[3] SHARE VSSI NCH L=60N W=1.5U M=4
MM17 YOUT[3] MWL2[3] VSSI VSSI NCH L=60N W=1.5U M=4
MM1 YOUT[2] PD_BUF VSSI VSSI NCH L=60N W=150.0N M=4
MM2 YOUT[3] PD_BUF VSSI VSSI NCH L=60N W=150.0N M=4
MM0 YOUT[1] PD_BUF VSSI VSSI NCH L=60N W=150.0N M=4
MN0 MWL2[0] YIN[0] SHARE VSSI NCH L=60N W=1.5U M=4
MN21 SHARE WLPY VSSI VSSI NCH L=60N W=600N M=16
MN19 YOUT[0] MWL2[0] VSSI VSSI NCH L=60N W=1.5U M=4
MN3 YOUT[0] PD_BUF VSSI VSSI NCH L=60N W=150.0N M=4
MM8 YOUT[2] MWL2[2] VSSI VSSI NCH L=60N W=1.5U M=4
MM7 YOUT[1] MWL2[1] VSSI VSSI NCH L=60N W=1.5U M=4
MM4 MWL2[1] YIN[1] SHARE VSSI NCH L=60N W=1.5U M=4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LCTRL
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LCTRL BLEQB_DN BLEQB_UP DEC_X3_DN DEC_X3_UP DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] 
+ DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] 
+ DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] 
+ DEC_Y_UP[6] DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLP_SAE 
+ YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO BLEQB_DN:I BLEQB_UP:I DEC_X3_DN:I DEC_X3_UP:I DEC_Y[0]:I DEC_Y[1]:I 
*.PININFO DEC_Y[2]:I DEC_Y[3]:I DEC_Y[4]:I DEC_Y[5]:I DEC_Y[6]:I DEC_Y[7]:I 
*.PININFO PD_BUF:I RW_RE:I WLP_SAE:I YL[0]:I DEC_Y_DN[0]:O DEC_Y_DN[1]:O 
*.PININFO DEC_Y_DN[2]:O DEC_Y_DN[3]:O DEC_Y_DN[4]:O DEC_Y_DN[5]:O 
*.PININFO DEC_Y_DN[6]:O DEC_Y_DN[7]:O DEC_Y_UP[0]:O DEC_Y_UP[1]:O 
*.PININFO DEC_Y_UP[2]:O DEC_Y_UP[3]:O DEC_Y_UP[4]:O DEC_Y_UP[5]:O 
*.PININFO DEC_Y_UP[6]:O DEC_Y_UP[7]:O RE:O SAEB:O WE:O YL_LIO[0]:O YL_LIO[1]:O 
*.PININFO VDDHD:B VDDI:B VSSI:B
XXDRV_READ BSD PD_BUF SAEB VDDHD VDDI VSSI WLP_SAE S1AHSF400W40_XDRV_READ
XXDRV_YL BS0 PD_BUF VDDHD VSSI YL[0] YL_LIO[0] YL_LIO[1] S1AHSF400W40_XDRV_Y10
XXDRV_RW BSD PD_BUF RE VDDHD VSSI WE RW_RE S1AHSF400W40_XDRV_RW
XXDRV_Y4_U<0> PD_BUF VDDHD VSSI BLEQB_UP DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] S1AHSF400W40_XDRV_Y4
XXDRV_Y4_U<1> PD_BUF VDDHD VSSI BLEQB_UP DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] 
+ DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] S1AHSF400W40_XDRV_Y4
XXDRV_Y4_D<0> PD_BUF VDDHD VSSI BLEQB_DN DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] S1AHSF400W40_XDRV_Y4
XXDRV_Y4_D<1> PD_BUF VDDHD VSSI BLEQB_DN DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] S1AHSF400W40_XDRV_Y4
XI229 BS3B VSSI VDDHD BS4 S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.6U LP=0.06U 
+ M=1
XI227 BS1B VSSI VDDHD BS2 S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.6U LP=0.06U 
+ M=1
XI228 BS2 VSSI VDDHD BS3B S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.6U LP=0.06U 
+ M=1
XINV0 BS0 VSSI VDDHD BS1B S1AHSF400W40_AINV FN=1 WN=0.3U LN=0.06U FP=1 WP=0.6U LP=0.06U 
+ M=1
XNAND0 BS0 BS4 VSSI VDDHD BSD S1AHSF400W40_ANAND FN2=2 WN2=1.2U LN2=0.06U FN1=2 WN1=1.2U 
+ LN1=0.06U FP1=2 WP1=1.2U LP1=0.06U FP2=2 WP2=1.2U LP2=0.06U M=1
XNOR0 DEC_X3_UP DEC_X3_DN VSSI VDDHD BS0 S1AHSF400W40_ANOR FN2=1 WN2=1U LN2=0.06U FN1=1 
+ WN1=1U LN1=0.06U FP1=1 WP1=1.2U LP1=0.06U FP2=1 WP2=1.2U LP2=0.06U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LCTRL_F_M8
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LCTRL_F_M8 BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] 
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] 
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] 
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF PD_CVDDBUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] 
+ WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE 
+ WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO DEC_Y[0]:I DEC_Y[1]:I DEC_Y[2]:I DEC_Y[3]:I DEC_Y[4]:I DEC_Y[5]:I 
*.PININFO DEC_Y[6]:I DEC_Y[7]:I PD_CVDDBUF:I YL[0]:I BLEQ_DN:O BLEQ_UP:O 
*.PININFO DEC_Y_DN[0]:O DEC_Y_DN[1]:O DEC_Y_DN[2]:O DEC_Y_DN[3]:O 
*.PININFO DEC_Y_DN[4]:O DEC_Y_DN[5]:O DEC_Y_DN[6]:O DEC_Y_DN[7]:O 
*.PININFO DEC_Y_UP[0]:O DEC_Y_UP[1]:O DEC_Y_UP[2]:O DEC_Y_UP[3]:O 
*.PININFO DEC_Y_UP[4]:O DEC_Y_UP[5]:O DEC_Y_UP[6]:O DEC_Y_UP[7]:O RE:O SAEB:O 
*.PININFO WE:O WLPY_DN[0]:O WLPY_DN[1]:O WLPY_DN[2]:O WLPY_DN[3]:O 
*.PININFO WLPY_UP[0]:O WLPY_UP[1]:O WLPY_UP[2]:O WLPY_UP[3]:O YL_LIO[0]:O 
*.PININFO YL_LIO[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B PD_BUF:B RW_RE:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B
XXDRV_WLP_U BLEQ_UP BLEQB_UP DEC_X3[1] PD_BUF WLP_SAE VDDHD VDDI VSSI 
+ WLPY_UP[0] S1AHSF400W40_XDRV_WLP_F
XXDRV_WLP_D BLEQ_DN BLEQB_DN DEC_X3[0] PD_BUF WLP_SAE VDDHD VDDI VSSI 
+ WLPY_DN[0] S1AHSF400W40_XDRV_WLP_F
XLCNT BLEQB_DN BLEQB_UP DEC_X3[0] DEC_X3[1] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] 
+ DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] 
+ DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] 
+ DEC_Y_UP[6] DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLP_SAE 
+ YL[0] YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LCTRL_F_M16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LCTRL_F_M16 BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] 
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] 
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] 
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF PD_CVDDBUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] 
+ WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE 
+ WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO DEC_X2[0]:I DEC_X2[1]:I DEC_X2[2]:I DEC_X2[3]:I DEC_Y[0]:I 
*.PININFO DEC_Y[1]:I DEC_Y[2]:I DEC_Y[3]:I DEC_Y[4]:I DEC_Y[5]:I DEC_Y[6]:I 
*.PININFO DEC_Y[7]:I PD_BUF:I PD_CVDDBUF:I RW_RE:I WLP_SAE:I WLP_SAE_TK:I 
*.PININFO YL[0]:I BLEQ_DN:O BLEQ_UP:O DEC_Y_DN[0]:O DEC_Y_DN[1]:O 
*.PININFO DEC_Y_DN[2]:O DEC_Y_DN[3]:O DEC_Y_DN[4]:O DEC_Y_DN[5]:O 
*.PININFO DEC_Y_DN[6]:O DEC_Y_DN[7]:O DEC_Y_UP[0]:O DEC_Y_UP[1]:O 
*.PININFO DEC_Y_UP[2]:O DEC_Y_UP[3]:O DEC_Y_UP[4]:O DEC_Y_UP[5]:O 
*.PININFO DEC_Y_UP[6]:O DEC_Y_UP[7]:O RE:O SAEB:O WE:O WLPY_DN[0]:O 
*.PININFO WLPY_DN[1]:O WLPY_DN[2]:O WLPY_DN[3]:O WLPY_UP[0]:O WLPY_UP[1]:O 
*.PININFO WLPY_UP[2]:O WLPY_UP[3]:O YL_LIO[0]:O YL_LIO[1]:O DEC_X0[0]:B 
*.PININFO DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B DEC_X0[5]:B 
*.PININFO DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B DEC_X1[2]:B 
*.PININFO DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B DEC_X1[7]:B 
*.PININFO DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B DEC_X3[4]:B 
*.PININFO DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B VDDHD:B VDDI:B VSSI:B
XLCTRL_F_M8 BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] 
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF PD_CVDDBUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] 
+ WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE 
+ WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL_F_M8
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_LCNT_M16_S64_D
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_LCNT_M16_S64_D BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] 
+ DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] 
+ DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] 
+ DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPYB_DN WLPYB_UP 
+ WLPY_DN WLPY_UP WLP_SAE WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO BLEQ_DN:B BLEQ_UP:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B DEC_Y_DN[0]:B DEC_Y_DN[1]:B DEC_Y_DN[2]:B DEC_Y_DN[3]:B 
*.PININFO DEC_Y_DN[4]:B DEC_Y_DN[5]:B DEC_Y_DN[6]:B DEC_Y_DN[7]:B 
*.PININFO DEC_Y_UP[0]:B DEC_Y_UP[1]:B DEC_Y_UP[2]:B DEC_Y_UP[3]:B 
*.PININFO DEC_Y_UP[4]:B DEC_Y_UP[5]:B DEC_Y_UP[6]:B DEC_Y_UP[7]:B PD_BUF:B 
*.PININFO RE:B RW_RE:B SAEB:B VDDHD:B VDDI:B VSSI:B WE:B WLPYB_DN:B WLPYB_UP:B 
*.PININFO WLPY_DN:B WLPY_UP:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B YL_LIO[0]:B 
*.PININFO YL_LIO[1]:B
XLCNT BLEQ_DN BLEQ_UP NET049[0] NET049[1] NET049[2] NET049[3] NET049[4] 
+ NET049[5] NET049[6] NET049[7] NET048[0] NET048[1] NET048[2] NET048[3] 
+ NET048[4] NET048[5] NET048[6] NET048[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] NET045[0] NET045[1] NET045[2] NET045[3] 
+ NET045[4] NET045[5] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF NET46 RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN WLPY_1[1] WLPY_1[2] 
+ WLPY_1[3] WLPY_UP WLPY_2[1] WLPY_2[2] WLPY_2[3] WLP_SAE NET010 YL[0] 
+ YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL_F_M16
XI3 VDDHD VDDI VSSI WLPY_UP WLPYB_UP S1AHSF400W40_XDRV_STRAP
XXDRV_STRP VDDHD VDDI VSSI WLPY_DN WLPYB_DN S1AHSF400W40_XDRV_STRAP
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_LCNT_M8_S64_D
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_LCNT_M8_S64_D BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] 
+ DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] 
+ DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] 
+ DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPYB_DN WLPYB_UP 
+ WLPY_DN WLPY_UP WLP_SAE WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO BLEQ_DN:B BLEQ_UP:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B DEC_Y_DN[0]:B DEC_Y_DN[1]:B DEC_Y_DN[2]:B DEC_Y_DN[3]:B 
*.PININFO DEC_Y_DN[4]:B DEC_Y_DN[5]:B DEC_Y_DN[6]:B DEC_Y_DN[7]:B 
*.PININFO DEC_Y_UP[0]:B DEC_Y_UP[1]:B DEC_Y_UP[2]:B DEC_Y_UP[3]:B 
*.PININFO DEC_Y_UP[4]:B DEC_Y_UP[5]:B DEC_Y_UP[6]:B DEC_Y_UP[7]:B PD_BUF:B 
*.PININFO RE:B RW_RE:B SAEB:B VDDHD:B VDDI:B VSSI:B WE:B WLPYB_DN:B WLPYB_UP:B 
*.PININFO WLPY_DN:B WLPY_UP:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B YL_LIO[0]:B 
*.PININFO YL_LIO[1]:B
XLCNT BLEQ_DN BLEQ_UP NET049[0] NET049[1] NET049[2] NET049[3] NET049[4] 
+ NET049[5] NET049[6] NET049[7] NET048[0] NET048[1] NET048[2] NET048[3] 
+ NET048[4] NET048[5] NET048[6] NET048[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] NET046[0] NET046[1] NET046[2] NET046[3] 
+ NET046[4] NET046[5] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF NET45 RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN WLPY_1[1] WLPY_1[2] 
+ WLPY_1[3] WLPY_UP WLPY_2[1] WLPY_2[2] WLPY_2[3] WLP_SAE NET045 YL[0] 
+ YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL_F_M8
XI3 VDDHD VDDI VSSI WLPY_UP WLPYB_UP S1AHSF400W40_XDRV_STRAP
XXDRV_STRP VDDHD VDDI VSSI WLPY_DN WLPYB_DN S1AHSF400W40_XDRV_STRAP
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LCTRL_F_M4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LCTRL_F_M4 BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] 
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] 
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] 
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF PD_CVDDBUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] 
+ WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE 
+ WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO DEC_Y[0]:I DEC_Y[1]:I DEC_Y[2]:I DEC_Y[3]:I DEC_Y[4]:I DEC_Y[5]:I 
*.PININFO DEC_Y[6]:I DEC_Y[7]:I PD_CVDDBUF:I YL[0]:I BLEQ_DN:O BLEQ_UP:O 
*.PININFO DEC_Y_DN[0]:O DEC_Y_DN[1]:O DEC_Y_DN[2]:O DEC_Y_DN[3]:O 
*.PININFO DEC_Y_DN[4]:O DEC_Y_DN[5]:O DEC_Y_DN[6]:O DEC_Y_DN[7]:O 
*.PININFO DEC_Y_UP[0]:O DEC_Y_UP[1]:O DEC_Y_UP[2]:O DEC_Y_UP[3]:O 
*.PININFO DEC_Y_UP[4]:O DEC_Y_UP[5]:O DEC_Y_UP[6]:O DEC_Y_UP[7]:O RE:O SAEB:O 
*.PININFO WE:O WLPY_DN[0]:O WLPY_DN[1]:O WLPY_DN[2]:O WLPY_DN[3]:O 
*.PININFO WLPY_UP[0]:O WLPY_UP[1]:O WLPY_UP[2]:O WLPY_UP[3]:O YL_LIO[0]:O 
*.PININFO YL_LIO[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B PD_BUF:B RW_RE:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B
XLCNT BLEQB_DN BLEQB_UP DEC_X3[0] DEC_X3[1] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] 
+ DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] 
+ DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] 
+ DEC_Y_UP[6] DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLP_SAE 
+ YL[0] YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL
XXDRV_WLP_U BLEQ_UP BLEQB_UP DEC_X3[1] PD_BUF WLP_SAE VDDHD VDDI VSSI 
+ WLPY_UP[0] S1AHSF400W40_XDRV_WLP_F
XXDRV_WLP_D BLEQ_DN BLEQB_DN DEC_X3[0] PD_BUF WLP_SAE VDDHD VDDI VSSI 
+ WLPY_DN[0] S1AHSF400W40_XDRV_WLP_F
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_LCNT_M4_S64_D
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_LCNT_M4_S64_D BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] 
+ DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] 
+ DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] 
+ DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPYB_DN WLPYB_UP 
+ WLPY_DN WLPY_UP WLP_SAE WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO BLEQ_DN:B BLEQ_UP:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B DEC_Y_DN[0]:B DEC_Y_DN[1]:B DEC_Y_DN[2]:B DEC_Y_DN[3]:B 
*.PININFO DEC_Y_DN[4]:B DEC_Y_DN[5]:B DEC_Y_DN[6]:B DEC_Y_DN[7]:B 
*.PININFO DEC_Y_UP[0]:B DEC_Y_UP[1]:B DEC_Y_UP[2]:B DEC_Y_UP[3]:B 
*.PININFO DEC_Y_UP[4]:B DEC_Y_UP[5]:B DEC_Y_UP[6]:B DEC_Y_UP[7]:B PD_BUF:B 
*.PININFO RE:B RW_RE:B SAEB:B VDDHD:B VDDI:B VSSI:B WE:B WLPYB_DN:B WLPYB_UP:B 
*.PININFO WLPY_DN:B WLPY_UP:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B YL_LIO[0]:B 
*.PININFO YL_LIO[1]:B
XLCNT BLEQ_DN BLEQ_UP NET049[0] NET049[1] NET049[2] NET049[3] NET049[4] 
+ NET049[5] NET049[6] NET049[7] NET048[0] NET048[1] NET048[2] NET048[3] 
+ NET048[4] NET048[5] NET048[6] NET048[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] NET046[0] NET046[1] NET046[2] NET046[3] 
+ NET046[4] NET046[5] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF NET45 RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN WLPY_1[1] WLPY_1[2] 
+ WLPY_1[3] WLPY_UP WLPY_2[1] WLPY_2[2] WLPY_2[3] WLP_SAE NET045 YL[0] 
+ YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL_F_M4
XI3 VDDHD VDDI VSSI WLPY_UP WLPYB_UP S1AHSF400W40_XDRV_STRAP
XXDRV_STRP VDDHD VDDI VSSI WLPY_DN WLPYB_DN S1AHSF400W40_XDRV_STRAP
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    XDRV_WLP_S
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_XDRV_WLP_S BLEQ BLEQB BS DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ PD_BUF RD_RST VDDHD VDDI VSSI WLOUT[0] WLOUT[1] WLOUT[2] WLOUT[3]
*.PININFO BS:I DEC_X2[0]:I DEC_X2[1]:I DEC_X2[2]:I DEC_X2[3]:I PD_BUF:I 
*.PININFO RD_RST:I BLEQ:O BLEQB:O WLOUT[0]:O WLOUT[1]:O WLOUT[2]:O WLOUT[3]:O 
*.PININFO VDDHD:B VDDI:B VSSI:B
MM4 MWL2[3] DEC_X2[3] VDDHD VDDHD PCH L=60N W=750.0N M=4
MM11 WLOUT[1] MWL2[1] VDDHD VDDHD PCH L=60N W=3U M=4
MM7 VDDHD RD_RSTB MWL2[2] VDDHD PCH L=60N W=750.0N M=4
MP20 BLEQB NET170 VDDHD VDDHD PCH L=60N W=750.0N M=8
MM3 MWL2[2] DEC_X2[2] VDDHD VDDHD PCH L=60N W=750.0N M=4
MM15 WLOUT[3] MWL2[3] VDDHD VDDHD PCH L=60N W=3U M=4
MM8 VDDHD RD_RSTB MWL2[3] VDDHD PCH L=60N W=750.0N M=4
MM14 WLOUT[2] MWL2[2] VDDHD VDDHD PCH L=60N W=3U M=4
MP21 BLEQB BSB VDDHD VDDHD PCH L=60N W=750.0N M=8
MM6 VDDHD RD_RSTB MWL2[1] VDDHD PCH L=60N W=750.0N M=4
MP28 WLOUT[0] MWL2[0] VDDHD VDDHD PCH L=60N W=3U M=4
MP16 MWL2[0] DEC_X2[0] VDDHD VDDHD PCH L=60N W=750.0N M=4
MP30 VDDHD RD_RSTB MWL2[0] VDDHD PCH L=60N W=750.0N M=4
MP31 SHARE RD_RSTB VDDHD VDDHD PCH L=60N W=750.0N M=1
MM0 MWL2[1] DEC_X2[1] VDDHD VDDHD PCH L=60N W=750.0N M=4
MM5 MWL2[3] DEC_X2[3] SHARE VSSI NCH L=60N W=1.5U M=4
MM13 WLOUT[2] MWL2[2] VSSI VSSI NCH L=60N W=1.5U M=4
MM12 WLOUT[1] MWL2[1] VSSI VSSI NCH L=60N W=1.5U M=4
MM16 WLOUT[3] MWL2[3] VSSI VSSI NCH L=60N W=1.5U M=4
MN21 SHARE RD_RSTB VSSI VSSI NCH L=60N W=600N M=16
MN19 WLOUT[0] MWL2[0] VSSI VSSI NCH L=60N W=1.5U M=4
MM1 MWL2[1] DEC_X2[1] SHARE VSSI NCH L=60N W=1.5U M=4
MN0 MWL2[0] DEC_X2[0] SHARE VSSI NCH L=60N W=1.5U M=4
MM2 MWL2[2] DEC_X2[2] SHARE VSSI NCH L=60N W=1.5U M=4
MN18 BLEQB BSB NET185 VSSI NCH L=60N W=750.0N M=8
MN2 NET185 NET170 VSSI VSSI NCH L=60N W=750.0N M=8
MN22 BLEQB PD_BUF VSSI VSSI NCH L=60N W=300N M=1
XI528 BS VSSI VDDHD BSB S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U LP=0.06U M=2
XINV2 BLEQB VSSI VDDI BLEQ S1AHSF400W40_AINV FN=8 WN=1.6U LN=0.07U FP=15 WP=1.6U LP=0.07U 
+ M=1
XINV1 NET149 VSSI VDDHD NET170 S1AHSF400W40_AINV FN=1 WN=1.2U LN=0.06U FP=1 WP=2.4U 
+ LP=0.06U M=1
XNAND0 NET160 NET156 VSSI VDDHD NET149 S1AHSF400W40_ANAND FN2=1 WN2=0.6U LN2=0.06U FN1=1 
+ WN1=0.6U LN1=0.06U FP1=1 WP1=1.2U LP1=0.06U FP2=1 WP2=1.2U LP2=0.06U M=1
XI527 BSB RD_RST VSSI VDDHD RD_RSTB S1AHSF400W40_ANOR FN2=2 WN2=0.5U LN2=0.06U FN1=2 
+ WN1=0.5U LN1=0.06U FP1=2 WP1=1.5U LP1=0.06U FP2=2 WP2=1.5U LP2=0.06U M=1
XI530 WLOUT[1] WLOUT[0] VSSI VDDHD NET156 S1AHSF400W40_ANOR FN2=1 WN2=0.3U LN2=0.06U 
+ FN1=1 WN1=0.3U LN1=0.06U FP1=1 WP1=1.2U LP1=0.06U FP2=1 WP2=1.2U LP2=0.06U 
+ M=1
XNOR1 WLOUT[2] WLOUT[3] VSSI VDDHD NET160 S1AHSF400W40_ANOR FN2=1 WN2=0.3U LN2=0.06U 
+ FN1=1 WN1=0.3U LN1=0.06U FP1=1 WP1=1.2U LP1=0.06U FP2=1 WP2=1.2U LP2=0.06U 
+ M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LCTRL_S_M8
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LCTRL_S_M8 BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] 
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] 
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] 
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF PD_CVDDBUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] 
+ WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE 
+ WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO DEC_Y[0]:I DEC_Y[1]:I DEC_Y[2]:I DEC_Y[3]:I DEC_Y[4]:I DEC_Y[5]:I 
*.PININFO DEC_Y[6]:I DEC_Y[7]:I PD_CVDDBUF:I YL[0]:I BLEQ_DN:O BLEQ_UP:O 
*.PININFO DEC_Y_DN[0]:O DEC_Y_DN[1]:O DEC_Y_DN[2]:O DEC_Y_DN[3]:O 
*.PININFO DEC_Y_DN[4]:O DEC_Y_DN[5]:O DEC_Y_DN[6]:O DEC_Y_DN[7]:O 
*.PININFO DEC_Y_UP[0]:O DEC_Y_UP[1]:O DEC_Y_UP[2]:O DEC_Y_UP[3]:O 
*.PININFO DEC_Y_UP[4]:O DEC_Y_UP[5]:O DEC_Y_UP[6]:O DEC_Y_UP[7]:O RE:O SAEB:O 
*.PININFO WE:O WLPY_DN[0]:O WLPY_DN[1]:O WLPY_DN[2]:O WLPY_DN[3]:O 
*.PININFO WLPY_UP[0]:O WLPY_UP[1]:O WLPY_UP[2]:O WLPY_UP[3]:O YL_LIO[0]:O 
*.PININFO YL_LIO[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B PD_BUF:B RW_RE:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B
XXDRV_WLP_UP BLEQ_UP BLEQB_UP DEC_X3[1] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] PD_BUF WLP_SAE VDDHD VDDI VSSI WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] 
+ WLPY_UP[3] S1AHSF400W40_XDRV_WLP_S
XXDRV_WLP_DN BLEQ_DN BLEQB_DN DEC_X3[0] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] PD_BUF WLP_SAE VDDHD VDDI VSSI WLPY_DN[0] WLPY_DN[1] WLPY_DN[2] 
+ WLPY_DN[3] S1AHSF400W40_XDRV_WLP_S
XLCTRL BLEQB_DN BLEQB_UP DEC_X3[0] DEC_X3[1] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] 
+ DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] 
+ DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] 
+ DEC_Y_UP[6] DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLP_SAE 
+ YL[0] YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_LCNT_M8_S256_D
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_LCNT_M8_S256_D BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] 
+ DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] 
+ DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] 
+ DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPYB_DN WLPYB_UP 
+ WLPY_DN WLPY_UP WLP_SAE WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO BLEQ_DN:B BLEQ_UP:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B DEC_Y_DN[0]:B DEC_Y_DN[1]:B DEC_Y_DN[2]:B DEC_Y_DN[3]:B 
*.PININFO DEC_Y_DN[4]:B DEC_Y_DN[5]:B DEC_Y_DN[6]:B DEC_Y_DN[7]:B 
*.PININFO DEC_Y_UP[0]:B DEC_Y_UP[1]:B DEC_Y_UP[2]:B DEC_Y_UP[3]:B 
*.PININFO DEC_Y_UP[4]:B DEC_Y_UP[5]:B DEC_Y_UP[6]:B DEC_Y_UP[7]:B PD_BUF:B 
*.PININFO RE:B RW_RE:B SAEB:B VDDHD:B VDDI:B VSSI:B WE:B WLPYB_DN:B WLPYB_UP:B 
*.PININFO WLPY_DN:B WLPY_UP:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B YL_LIO[0]:B 
*.PININFO YL_LIO[1]:B
XLCNT BLEQ_DN BLEQ_UP NET045[0] NET045[1] NET045[2] NET045[3] NET045[4] 
+ NET045[5] NET045[6] NET045[7] NET046[0] NET046[1] NET046[2] NET046[3] 
+ NET046[4] NET046[5] NET046[6] NET046[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] NET049[0] NET049[1] NET049[2] NET049[3] 
+ NET049[4] NET049[5] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF NET45 RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN WLPY_1[1] WLPY_1[2] 
+ WLPY_1[3] WLPY_2[0] WLPY_2[1] WLPY_2[2] WLPY_UP WLP_SAE NET010 YL[0] 
+ YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL_S_M8
XI3 VDDHD VDDI VSSI WLPY_UP WLPYB_UP S1AHSF400W40_XDRV_STRAP
XXDRV_STRP VDDHD VDDI VSSI WLPY_DN WLPYB_DN S1AHSF400W40_XDRV_STRAP
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LCTRL_S_M16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LCTRL_S_M16 BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] 
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] 
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] 
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF PD_CVDDBUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] 
+ WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE 
+ WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO DEC_X2[0]:I DEC_X2[1]:I DEC_X2[2]:I DEC_X2[3]:I DEC_Y[0]:I 
*.PININFO DEC_Y[1]:I DEC_Y[2]:I DEC_Y[3]:I DEC_Y[4]:I DEC_Y[5]:I DEC_Y[6]:I 
*.PININFO DEC_Y[7]:I PD_BUF:I PD_CVDDBUF:I RW_RE:I WLP_SAE:I WLP_SAE_TK:I 
*.PININFO YL[0]:I BLEQ_DN:O BLEQ_UP:O DEC_Y_DN[0]:O DEC_Y_DN[1]:O 
*.PININFO DEC_Y_DN[2]:O DEC_Y_DN[3]:O DEC_Y_DN[4]:O DEC_Y_DN[5]:O 
*.PININFO DEC_Y_DN[6]:O DEC_Y_DN[7]:O DEC_Y_UP[0]:O DEC_Y_UP[1]:O 
*.PININFO DEC_Y_UP[2]:O DEC_Y_UP[3]:O DEC_Y_UP[4]:O DEC_Y_UP[5]:O 
*.PININFO DEC_Y_UP[6]:O DEC_Y_UP[7]:O RE:O SAEB:O WE:O WLPY_DN[0]:O 
*.PININFO WLPY_DN[1]:O WLPY_DN[2]:O WLPY_DN[3]:O WLPY_UP[0]:O WLPY_UP[1]:O 
*.PININFO WLPY_UP[2]:O WLPY_UP[3]:O YL_LIO[0]:O YL_LIO[1]:O DEC_X0[0]:B 
*.PININFO DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B DEC_X0[5]:B 
*.PININFO DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B DEC_X1[2]:B 
*.PININFO DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B DEC_X1[7]:B 
*.PININFO DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B DEC_X3[4]:B 
*.PININFO DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B VDDHD:B VDDI:B VSSI:B
XLCTRL_S_M8 BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] 
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF PD_CVDDBUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] 
+ WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE 
+ WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL_S_M8
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_LCNT_M16_S256_D
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_LCNT_M16_S256_D BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] 
+ DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] 
+ DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] 
+ DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPYB_DN WLPYB_UP 
+ WLPY_DN WLPY_UP WLP_SAE WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO BLEQ_DN:B BLEQ_UP:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B DEC_Y_DN[0]:B DEC_Y_DN[1]:B DEC_Y_DN[2]:B DEC_Y_DN[3]:B 
*.PININFO DEC_Y_DN[4]:B DEC_Y_DN[5]:B DEC_Y_DN[6]:B DEC_Y_DN[7]:B 
*.PININFO DEC_Y_UP[0]:B DEC_Y_UP[1]:B DEC_Y_UP[2]:B DEC_Y_UP[3]:B 
*.PININFO DEC_Y_UP[4]:B DEC_Y_UP[5]:B DEC_Y_UP[6]:B DEC_Y_UP[7]:B PD_BUF:B 
*.PININFO RE:B RW_RE:B SAEB:B VDDHD:B VDDI:B VSSI:B WE:B WLPYB_DN:B WLPYB_UP:B 
*.PININFO WLPY_DN:B WLPY_UP:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B YL_LIO[0]:B 
*.PININFO YL_LIO[1]:B
XLCNT BLEQ_DN BLEQ_UP NET049[0] NET049[1] NET049[2] NET049[3] NET049[4] 
+ NET049[5] NET049[6] NET049[7] NET045[0] NET045[1] NET045[2] NET045[3] 
+ NET045[4] NET045[5] NET045[6] NET045[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] NET048[0] NET048[1] NET048[2] NET048[3] 
+ NET048[4] NET048[5] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF NET45 RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN WLPY_1[1] WLPY_1[2] 
+ WLPY_1[3] WLPY_2[0] WLPY_2[1] WLPY_2[2] WLPY_UP WLP_SAE NET010 YL[0] 
+ YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL_S_M16
XI3 VDDHD VDDI VSSI WLPY_UP WLPYB_UP S1AHSF400W40_XDRV_STRAP
XXDRV_STRP VDDHD VDDI VSSI WLPY_DN WLPYB_DN S1AHSF400W40_XDRV_STRAP
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LCTRL_S_M4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LCTRL_S_M4 BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] 
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] 
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] 
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF PD_CVDDBUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] 
+ WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE 
+ WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO DEC_Y[0]:I DEC_Y[1]:I DEC_Y[2]:I DEC_Y[3]:I DEC_Y[4]:I DEC_Y[5]:I 
*.PININFO DEC_Y[6]:I DEC_Y[7]:I PD_CVDDBUF:I YL[0]:I BLEQ_DN:O BLEQ_UP:O 
*.PININFO DEC_Y_DN[0]:O DEC_Y_DN[1]:O DEC_Y_DN[2]:O DEC_Y_DN[3]:O 
*.PININFO DEC_Y_DN[4]:O DEC_Y_DN[5]:O DEC_Y_DN[6]:O DEC_Y_DN[7]:O 
*.PININFO DEC_Y_UP[0]:O DEC_Y_UP[1]:O DEC_Y_UP[2]:O DEC_Y_UP[3]:O 
*.PININFO DEC_Y_UP[4]:O DEC_Y_UP[5]:O DEC_Y_UP[6]:O DEC_Y_UP[7]:O RE:O SAEB:O 
*.PININFO WE:O WLPY_DN[0]:O WLPY_DN[1]:O WLPY_DN[2]:O WLPY_DN[3]:O 
*.PININFO WLPY_UP[0]:O WLPY_UP[1]:O WLPY_UP[2]:O WLPY_UP[3]:O YL_LIO[0]:O 
*.PININFO YL_LIO[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B PD_BUF:B RW_RE:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B
XLCTRL BLEQB_DN BLEQB_UP DEC_X3[0] DEC_X3[1] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] 
+ DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] 
+ DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] 
+ DEC_Y_UP[6] DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLP_SAE 
+ YL[0] YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL
XXDRV_WLP_UP BLEQ_UP BLEQB_UP DEC_X3[1] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] PD_BUF WLP_SAE VDDHD VDDI VSSI WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] 
+ WLPY_UP[3] S1AHSF400W40_XDRV_WLP_S
XXDRV_WLP_DN BLEQ_DN BLEQB_DN DEC_X3[0] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] PD_BUF WLP_SAE VDDHD VDDI VSSI WLPY_DN[0] WLPY_DN[1] WLPY_DN[2] 
+ WLPY_DN[3] S1AHSF400W40_XDRV_WLP_S
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_LCNT_M4_S256_D
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_LCNT_M4_S256_D BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] 
+ DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] 
+ DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] 
+ DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPYB_DN WLPYB_UP 
+ WLPY_DN WLPY_UP WLP_SAE WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO BLEQ_DN:B BLEQ_UP:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B DEC_Y_DN[0]:B DEC_Y_DN[1]:B DEC_Y_DN[2]:B DEC_Y_DN[3]:B 
*.PININFO DEC_Y_DN[4]:B DEC_Y_DN[5]:B DEC_Y_DN[6]:B DEC_Y_DN[7]:B 
*.PININFO DEC_Y_UP[0]:B DEC_Y_UP[1]:B DEC_Y_UP[2]:B DEC_Y_UP[3]:B 
*.PININFO DEC_Y_UP[4]:B DEC_Y_UP[5]:B DEC_Y_UP[6]:B DEC_Y_UP[7]:B PD_BUF:B 
*.PININFO RE:B RW_RE:B SAEB:B VDDHD:B VDDI:B VSSI:B WE:B WLPYB_DN:B WLPYB_UP:B 
*.PININFO WLPY_DN:B WLPY_UP:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B YL_LIO[0]:B 
*.PININFO YL_LIO[1]:B
XI3 VDDHD VDDI VSSI WLPY_UP WLPYB_UP S1AHSF400W40_XDRV_STRAP
XXDRV_STRP VDDHD VDDI VSSI WLPY_DN WLPYB_DN S1AHSF400W40_XDRV_STRAP
XLCNT BLEQ_DN BLEQ_UP NET060[0] NET060[1] NET060[2] NET060[3] NET060[4] 
+ NET060[5] NET060[6] NET060[7] NET061[0] NET061[1] NET061[2] NET061[3] 
+ NET061[4] NET061[5] NET061[6] NET061[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] NET059[0] NET059[1] NET059[2] NET059[3] 
+ NET059[4] NET059[5] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF NET45 RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN WLPY_1[1] WLPY_1[2] 
+ WLPY_1[3] WLPY_2[0] WLPY_2[1] WLPY_2[2] WLPY_UP WLP_SAE NET057 YL[0] 
+ YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL_S_M4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_LCNT_D_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_LCNT_D_SIM BLEQ_DN_LT BLEQ_DN_RT BLEQ_UP_LT BLEQ_UP_RT CVDDHD CVDDI 
+ DEC_X0_BT[0] DEC_X0_BT[1] DEC_X0_BT[2] DEC_X0_BT[3] DEC_X0_BT[4] 
+ DEC_X0_BT[5] DEC_X0_BT[6] DEC_X0_BT[7] DEC_X0_TP[0] DEC_X0_TP[1] 
+ DEC_X0_TP[2] DEC_X0_TP[3] DEC_X0_TP[4] DEC_X0_TP[5] DEC_X0_TP[6] 
+ DEC_X0_TP[7] DEC_X1_BT[0] DEC_X1_BT[1] DEC_X1_BT[2] DEC_X1_BT[3] 
+ DEC_X1_BT[4] DEC_X1_BT[5] DEC_X1_BT[6] DEC_X1_BT[7] DEC_X1_TP[0] 
+ DEC_X1_TP[1] DEC_X1_TP[2] DEC_X1_TP[3] DEC_X1_TP[4] DEC_X1_TP[5] 
+ DEC_X1_TP[6] DEC_X1_TP[7] DEC_X2_BT[0] DEC_X2_BT[1] DEC_X2_BT[2] 
+ DEC_X2_BT[3] DEC_X2_TP[0] DEC_X2_TP[1] DEC_X2_TP[2] DEC_X2_TP[3] 
+ DEC_X3_BT[0] DEC_X3_BT[1] DEC_X3_BT[2] DEC_X3_BT[3] DEC_X3_BT[4] 
+ DEC_X3_BT[5] DEC_X3_BT[6] DEC_X3_BT[7] DEC_X3_TP[0] DEC_X3_TP[1] 
+ DEC_X3_TP[2] DEC_X3_TP[3] DEC_X3_TP[4] DEC_X3_TP[5] DEC_X3_TP[6] 
+ DEC_X3_TP[7] DEC_Y_BT[0] DEC_Y_BT[1] DEC_Y_BT[2] DEC_Y_BT[3] DEC_Y_BT[4] 
+ DEC_Y_BT[5] DEC_Y_BT[6] DEC_Y_BT[7] DEC_Y_DN_LT[0] DEC_Y_DN_LT[1] 
+ DEC_Y_DN_LT[2] DEC_Y_DN_LT[3] DEC_Y_DN_LT[4] DEC_Y_DN_LT[5] DEC_Y_DN_LT[6] 
+ DEC_Y_DN_LT[7] DEC_Y_DN_RT[0] DEC_Y_DN_RT[1] DEC_Y_DN_RT[2] DEC_Y_DN_RT[3] 
+ DEC_Y_DN_RT[4] DEC_Y_DN_RT[5] DEC_Y_DN_RT[6] DEC_Y_DN_RT[7] DEC_Y_TP[0] 
+ DEC_Y_TP[1] DEC_Y_TP[2] DEC_Y_TP[3] DEC_Y_TP[4] DEC_Y_TP[5] DEC_Y_TP[6] 
+ DEC_Y_TP[7] DEC_Y_UP_LT[0] DEC_Y_UP_LT[1] DEC_Y_UP_LT[2] DEC_Y_UP_LT[3] 
+ DEC_Y_UP_LT[4] DEC_Y_UP_LT[5] DEC_Y_UP_LT[6] DEC_Y_UP_LT[7] DEC_Y_UP_RT[0] 
+ DEC_Y_UP_RT[1] DEC_Y_UP_RT[2] DEC_Y_UP_RT[3] DEC_Y_UP_RT[4] DEC_Y_UP_RT[5] 
+ DEC_Y_UP_RT[6] DEC_Y_UP_RT[7] PD_BUF_BT PD_BUF_TP PD_CVDDBUF_BT 
+ PD_CVDDBUF_TP RE_LT RE_RT RW_RE_BT RW_RE_TP SAEB_LT SAEB_RT VDDHD VDDI VSSI 
+ WE_LT WE_RT WLPYB_DN_BT WLPYB_UP_TP WLPY_DN_BT WLPY_UP_TP WLP_SAE_BT 
+ WLP_SAE_TK_BT WLP_SAE_TK_TP WLP_SAE_TP YL_BT[0] YL_LIO_LT[0] YL_LIO_LT[1] 
+ YL_LIO_RT[0] YL_LIO_RT[1] YL_TP[0]
*.PININFO DEC_X0_BT[0]:I DEC_X0_BT[1]:I DEC_X0_BT[2]:I DEC_X0_BT[3]:I 
*.PININFO DEC_X0_BT[4]:I DEC_X0_BT[5]:I DEC_X0_BT[6]:I DEC_X0_BT[7]:I 
*.PININFO DEC_X1_BT[0]:I DEC_X1_BT[1]:I DEC_X1_BT[2]:I DEC_X1_BT[3]:I 
*.PININFO DEC_X1_BT[4]:I DEC_X1_BT[5]:I DEC_X1_BT[6]:I DEC_X1_BT[7]:I 
*.PININFO PD_BUF_BT:I PD_CVDDBUF_BT:I RW_RE_TP:I DEC_X0_TP[0]:O DEC_X0_TP[1]:O 
*.PININFO DEC_X0_TP[2]:O DEC_X0_TP[3]:O DEC_X0_TP[4]:O DEC_X0_TP[5]:O 
*.PININFO DEC_X0_TP[6]:O DEC_X0_TP[7]:O DEC_X1_TP[0]:O DEC_X1_TP[1]:O 
*.PININFO DEC_X1_TP[2]:O DEC_X1_TP[3]:O DEC_X1_TP[4]:O DEC_X1_TP[5]:O 
*.PININFO DEC_X1_TP[6]:O DEC_X1_TP[7]:O PD_BUF_TP:O PD_CVDDBUF_TP:O 
*.PININFO BLEQ_DN_LT:B BLEQ_DN_RT:B BLEQ_UP_LT:B BLEQ_UP_RT:B CVDDHD:B CVDDI:B 
*.PININFO DEC_X2_BT[0]:B DEC_X2_BT[1]:B DEC_X2_BT[2]:B DEC_X2_BT[3]:B 
*.PININFO DEC_X2_TP[0]:B DEC_X2_TP[1]:B DEC_X2_TP[2]:B DEC_X2_TP[3]:B 
*.PININFO DEC_X3_BT[0]:B DEC_X3_BT[1]:B DEC_X3_BT[2]:B DEC_X3_BT[3]:B 
*.PININFO DEC_X3_BT[4]:B DEC_X3_BT[5]:B DEC_X3_BT[6]:B DEC_X3_BT[7]:B 
*.PININFO DEC_X3_TP[0]:B DEC_X3_TP[1]:B DEC_X3_TP[2]:B DEC_X3_TP[3]:B 
*.PININFO DEC_X3_TP[4]:B DEC_X3_TP[5]:B DEC_X3_TP[6]:B DEC_X3_TP[7]:B 
*.PININFO DEC_Y_BT[0]:B DEC_Y_BT[1]:B DEC_Y_BT[2]:B DEC_Y_BT[3]:B 
*.PININFO DEC_Y_BT[4]:B DEC_Y_BT[5]:B DEC_Y_BT[6]:B DEC_Y_BT[7]:B 
*.PININFO DEC_Y_DN_LT[0]:B DEC_Y_DN_LT[1]:B DEC_Y_DN_LT[2]:B DEC_Y_DN_LT[3]:B 
*.PININFO DEC_Y_DN_LT[4]:B DEC_Y_DN_LT[5]:B DEC_Y_DN_LT[6]:B DEC_Y_DN_LT[7]:B 
*.PININFO DEC_Y_DN_RT[0]:B DEC_Y_DN_RT[1]:B DEC_Y_DN_RT[2]:B DEC_Y_DN_RT[3]:B 
*.PININFO DEC_Y_DN_RT[4]:B DEC_Y_DN_RT[5]:B DEC_Y_DN_RT[6]:B DEC_Y_DN_RT[7]:B 
*.PININFO DEC_Y_TP[0]:B DEC_Y_TP[1]:B DEC_Y_TP[2]:B DEC_Y_TP[3]:B 
*.PININFO DEC_Y_TP[4]:B DEC_Y_TP[5]:B DEC_Y_TP[6]:B DEC_Y_TP[7]:B 
*.PININFO DEC_Y_UP_LT[0]:B DEC_Y_UP_LT[1]:B DEC_Y_UP_LT[2]:B DEC_Y_UP_LT[3]:B 
*.PININFO DEC_Y_UP_LT[4]:B DEC_Y_UP_LT[5]:B DEC_Y_UP_LT[6]:B DEC_Y_UP_LT[7]:B 
*.PININFO DEC_Y_UP_RT[0]:B DEC_Y_UP_RT[1]:B DEC_Y_UP_RT[2]:B DEC_Y_UP_RT[3]:B 
*.PININFO DEC_Y_UP_RT[4]:B DEC_Y_UP_RT[5]:B DEC_Y_UP_RT[6]:B DEC_Y_UP_RT[7]:B 
*.PININFO RE_LT:B RE_RT:B RW_RE_BT:B SAEB_LT:B SAEB_RT:B VDDHD:B VDDI:B VSSI:B 
*.PININFO WE_LT:B WE_RT:B WLPYB_DN_BT:B WLPYB_UP_TP:B WLPY_DN_BT:B 
*.PININFO WLPY_UP_TP:B WLP_SAE_BT:B WLP_SAE_TK_BT:B WLP_SAE_TK_TP:B 
*.PININFO WLP_SAE_TP:B YL_BT[0]:B YL_LIO_LT[0]:B YL_LIO_LT[1]:B YL_LIO_RT[0]:B 
*.PININFO YL_LIO_RT[1]:B YL_TP[0]:B
XI27 NET0181 NET0180 NET0179[0] NET0179[1] NET0179[2] NET0179[3] NET0179[4] 
+ NET0179[5] NET0179[6] NET0179[7] NET0178[0] NET0178[1] NET0178[2] NET0178[3] 
+ NET0178[4] NET0178[5] NET0178[6] NET0178[7] NET0177[0] NET0177[1] NET0177[2] 
+ NET0177[3] NET0176[0] NET0176[1] NET0176[2] NET0176[3] NET0176[4] NET0176[5] 
+ NET0176[6] NET0176[7] NET0175[0] NET0175[1] NET0175[2] NET0175[3] NET0175[4] 
+ NET0175[5] NET0175[6] NET0175[7] NET0174[0] NET0174[1] NET0174[2] NET0174[3] 
+ NET0174[4] NET0174[5] NET0174[6] NET0174[7] NET0173[0] NET0173[1] NET0173[2] 
+ NET0173[3] NET0173[4] NET0173[5] NET0173[6] NET0173[7] NET0172 NET0171 
+ NET0170 NET0169 NET0168 NET0167 NET0166 NET0182 NET0185 NET0184 NET0165 
+ NET0164 NET0163 NET0162 NET0161 NET0183[0] NET0183[1] S1AHSF400W40_BK_LCNT_M16_S64_D
XI26 NET081 NET080 NET079[0] NET079[1] NET079[2] NET079[3] NET079[4] NET079[5] 
+ NET079[6] NET079[7] NET078[0] NET078[1] NET078[2] NET078[3] NET078[4] 
+ NET078[5] NET078[6] NET078[7] NET011[0] NET011[1] NET011[2] NET011[3] 
+ NET076[0] NET076[1] NET076[2] NET076[3] NET076[4] NET076[5] NET076[6] 
+ NET076[7] NET075[0] NET075[1] NET075[2] NET075[3] NET075[4] NET075[5] 
+ NET075[6] NET075[7] NET074[0] NET074[1] NET074[2] NET074[3] NET074[4] 
+ NET074[5] NET074[6] NET074[7] NET073[0] NET073[1] NET073[2] NET073[3] 
+ NET073[4] NET073[5] NET073[6] NET073[7] NET072 NET09 NET018 NET019 NET014 
+ NET08 NET017 NET082 NET016 NET084 NET013 NET06 NET03 NET07 NET015 NET083[0] 
+ NET083[1] S1AHSF400W40_BK_LCNT_M8_S64_D
XI25 NET0106 NET0105 NET0104[0] NET0104[1] NET0104[2] NET0104[3] NET0104[4] 
+ NET0104[5] NET0104[6] NET0104[7] NET0103[0] NET0103[1] NET0103[2] NET0103[3] 
+ NET0103[4] NET0103[5] NET0103[6] NET0103[7] NET0102[0] NET0102[1] NET0102[2] 
+ NET0102[3] NET0101[0] NET0101[1] NET0101[2] NET0101[3] NET0101[4] NET0101[5] 
+ NET0101[6] NET0101[7] NET0100[0] NET0100[1] NET0100[2] NET0100[3] NET0100[4] 
+ NET0100[5] NET0100[6] NET0100[7] NET099[0] NET099[1] NET099[2] NET099[3] 
+ NET099[4] NET099[5] NET099[6] NET099[7] NET098[0] NET098[1] NET098[2] 
+ NET098[3] NET098[4] NET098[5] NET098[6] NET098[7] NET097 NET096 NET094 
+ NET093 NET092 NET091 NET090 NET0107 NET0110 NET0109 NET089 NET088 NET087 
+ NET095 NET086 NET0108[0] NET0108[1] S1AHSF400W40_BK_LCNT_M4_S64_D
XI24 NET0131 NET0130 NET0129[0] NET0129[1] NET0129[2] NET0129[3] NET0129[4] 
+ NET0129[5] NET0129[6] NET0129[7] NET0128[0] NET0128[1] NET0128[2] NET0128[3] 
+ NET0128[4] NET0128[5] NET0128[6] NET0128[7] NET0127[0] NET0127[1] NET0127[2] 
+ NET0127[3] NET0126[0] NET0126[1] NET0126[2] NET0126[3] NET0126[4] NET0126[5] 
+ NET0126[6] NET0126[7] NET0125[0] NET0125[1] NET0125[2] NET0125[3] NET0125[4] 
+ NET0125[5] NET0125[6] NET0125[7] NET0124[0] NET0124[1] NET0124[2] NET0124[3] 
+ NET0124[4] NET0124[5] NET0124[6] NET0124[7] NET0123[0] NET0123[1] NET0123[2] 
+ NET0123[3] NET0123[4] NET0123[5] NET0123[6] NET0123[7] NET0122 NET0121 
+ NET0120 NET0119 NET0118 NET0117 NET0116 NET0132 NET0135 NET0134 NET0115 
+ NET0114 NET0113 NET0112 NET0111 NET0133[0] NET0133[1] S1AHSF400W40_BK_LCNT_M8_S256_D
XI23 NET067 NET066 NET065[0] NET065[1] NET065[2] NET065[3] NET065[4] NET065[5] 
+ NET065[6] NET065[7] NET064[0] NET064[1] NET064[2] NET064[3] NET064[4] 
+ NET064[5] NET064[6] NET064[7] NET063[0] NET063[1] NET063[2] NET063[3] 
+ NET062[0] NET062[1] NET062[2] NET062[3] NET062[4] NET062[5] NET062[6] 
+ NET062[7] NET061[0] NET061[1] NET061[2] NET061[3] NET061[4] NET061[5] 
+ NET061[6] NET061[7] NET060[0] NET060[1] NET060[2] NET060[3] NET060[4] 
+ NET060[5] NET060[6] NET060[7] NET059[0] NET059[1] NET059[2] NET059[3] 
+ NET059[4] NET059[5] NET059[6] NET059[7] NET058 NET057 NET056 NET055 NET054 
+ NET053 NET052 NET068 NET071 NET070 NET051 NET04 NET05 NET010 NET012 
+ NET069[0] NET069[1] S1AHSF400W40_BK_LCNT_M16_S256_D
XI22 NET68 NET67 NET66[0] NET66[1] NET66[2] NET66[3] NET66[4] NET66[5] 
+ NET66[6] NET66[7] NET65[0] NET65[1] NET65[2] NET65[3] NET65[4] NET65[5] 
+ NET65[6] NET65[7] NET64[0] NET64[1] NET64[2] NET64[3] NET63[0] NET63[1] 
+ NET63[2] NET63[3] NET63[4] NET63[5] NET63[6] NET63[7] NET62[0] NET62[1] 
+ NET62[2] NET62[3] NET62[4] NET62[5] NET62[6] NET62[7] NET61[0] NET61[1] 
+ NET61[2] NET61[3] NET61[4] NET61[5] NET61[6] NET61[7] NET60[0] NET60[1] 
+ NET60[2] NET60[3] NET60[4] NET60[5] NET60[6] NET60[7] NET59 NET01 NET56 
+ NET55 NET54 NET53 NET52 NET02 NET049 NET048 NET047 NET046 NET48 NET085 
+ NET077 NET050[0] NET050[1] S1AHSF400W40_BK_LCNT_M4_S256_D
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    WLPY_32_LD
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_WLPY_32_LD VDDHD VDDI VSSI WLPYB_LD WLPY_LD
*.PININFO VDDHD:B VDDI:B VSSI:B WLPYB_LD:B WLPY_LD:B
XWLDV_0<0> NET05[0] NET018[0] NET017[0] NET017[1] NET017[2] NET017[3] 
+ NET017[4] NET017[5] NET04[0] NET015[0] NET015[1] NET015[2] NET015[3] 
+ NET015[4] NET015[5] NET015[6] NET011[0] NET011[1] NET011[2] NET011[3] 
+ NET012[0] NET012[1] NET012[2] NET012[3] NET012[4] NET012[5] NET012[6] 
+ NET012[7] NET014[0] NET014[1] NET014[2] NET014[3] NET014[4] NET014[5] 
+ NET014[6] NET014[7] NET03 NET016[0] NET010[0] VDDHD VDDI VSSI NET019[0] 
+ NET019[1] WLPY_LD WLPYB_LD NET09[0] NET07[0] NET013[0] S1AHSF400W40_XDRV_LA512
XWLDV_0<1> NET05[1] NET018[1] NET017[6] NET017[7] NET017[8] NET017[9] 
+ NET017[10] NET017[11] NET04[1] NET015[7] NET015[8] NET015[9] NET015[10] 
+ NET015[11] NET015[12] NET015[13] NET011[4] NET011[5] NET011[6] NET011[7] 
+ NET012[8] NET012[9] NET012[10] NET012[11] NET012[12] NET012[13] NET012[14] 
+ NET012[15] NET014[8] NET014[9] NET014[10] NET014[11] NET014[12] NET014[13] 
+ NET014[14] NET014[15] NET03 NET016[1] NET010[1] VDDHD VDDI VSSI NET019[2] 
+ NET019[3] WLPY_LD WLPYB_LD NET09[1] NET07[1] NET013[1] S1AHSF400W40_XDRV_LA512
XWLDV_0<2> NET05[2] NET018[2] NET017[12] NET017[13] NET017[14] NET017[15] 
+ NET017[16] NET017[17] NET04[2] NET015[14] NET015[15] NET015[16] NET015[17] 
+ NET015[18] NET015[19] NET015[20] NET011[8] NET011[9] NET011[10] NET011[11] 
+ NET012[16] NET012[17] NET012[18] NET012[19] NET012[20] NET012[21] NET012[22] 
+ NET012[23] NET014[16] NET014[17] NET014[18] NET014[19] NET014[20] NET014[21] 
+ NET014[22] NET014[23] NET03 NET016[2] NET010[2] VDDHD VDDI VSSI NET019[4] 
+ NET019[5] WLPY_LD WLPYB_LD NET09[2] NET07[2] NET013[2] S1AHSF400W40_XDRV_LA512
XWLDV_0<3> NET05[3] NET018[3] NET017[18] NET017[19] NET017[20] NET017[21] 
+ NET017[22] NET017[23] NET04[3] NET015[21] NET015[22] NET015[23] NET015[24] 
+ NET015[25] NET015[26] NET015[27] NET011[12] NET011[13] NET011[14] NET011[15] 
+ NET012[24] NET012[25] NET012[26] NET012[27] NET012[28] NET012[29] NET012[30] 
+ NET012[31] NET014[24] NET014[25] NET014[26] NET014[27] NET014[28] NET014[29] 
+ NET014[30] NET014[31] NET03 NET016[3] NET010[3] VDDHD VDDI VSSI NET019[6] 
+ NET019[7] WLPY_LD WLPYB_LD NET09[3] NET07[3] NET013[3] S1AHSF400W40_XDRV_LA512
XWLDV_0<4> NET05[4] NET018[4] NET017[24] NET017[25] NET017[26] NET017[27] 
+ NET017[28] NET017[29] NET04[4] NET015[28] NET015[29] NET015[30] NET015[31] 
+ NET015[32] NET015[33] NET015[34] NET011[16] NET011[17] NET011[18] NET011[19] 
+ NET012[32] NET012[33] NET012[34] NET012[35] NET012[36] NET012[37] NET012[38] 
+ NET012[39] NET014[32] NET014[33] NET014[34] NET014[35] NET014[36] NET014[37] 
+ NET014[38] NET014[39] NET03 NET016[4] NET010[4] VDDHD VDDI VSSI NET019[8] 
+ NET019[9] WLPY_LD WLPYB_LD NET09[4] NET07[4] NET013[4] S1AHSF400W40_XDRV_LA512
XWLDV_0<5> NET05[5] NET018[5] NET017[30] NET017[31] NET017[32] NET017[33] 
+ NET017[34] NET017[35] NET04[5] NET015[35] NET015[36] NET015[37] NET015[38] 
+ NET015[39] NET015[40] NET015[41] NET011[20] NET011[21] NET011[22] NET011[23] 
+ NET012[40] NET012[41] NET012[42] NET012[43] NET012[44] NET012[45] NET012[46] 
+ NET012[47] NET014[40] NET014[41] NET014[42] NET014[43] NET014[44] NET014[45] 
+ NET014[46] NET014[47] NET03 NET016[5] NET010[5] VDDHD VDDI VSSI NET019[10] 
+ NET019[11] WLPY_LD WLPYB_LD NET09[5] NET07[5] NET013[5] S1AHSF400W40_XDRV_LA512
XWLDV_0<6> NET05[6] NET018[6] NET017[36] NET017[37] NET017[38] NET017[39] 
+ NET017[40] NET017[41] NET04[6] NET015[42] NET015[43] NET015[44] NET015[45] 
+ NET015[46] NET015[47] NET015[48] NET011[24] NET011[25] NET011[26] NET011[27] 
+ NET012[48] NET012[49] NET012[50] NET012[51] NET012[52] NET012[53] NET012[54] 
+ NET012[55] NET014[48] NET014[49] NET014[50] NET014[51] NET014[52] NET014[53] 
+ NET014[54] NET014[55] NET03 NET016[6] NET010[6] VDDHD VDDI VSSI NET019[12] 
+ NET019[13] WLPY_LD WLPYB_LD NET09[6] NET07[6] NET013[6] S1AHSF400W40_XDRV_LA512
XWLDV_0<7> NET05[7] NET018[7] NET017[42] NET017[43] NET017[44] NET017[45] 
+ NET017[46] NET017[47] NET04[7] NET015[49] NET015[50] NET015[51] NET015[52] 
+ NET015[53] NET015[54] NET015[55] NET011[28] NET011[29] NET011[30] NET011[31] 
+ NET012[56] NET012[57] NET012[58] NET012[59] NET012[60] NET012[61] NET012[62] 
+ NET012[63] NET014[56] NET014[57] NET014[58] NET014[59] NET014[60] NET014[61] 
+ NET014[62] NET014[63] NET03 NET016[7] NET010[7] VDDHD VDDI VSSI NET019[14] 
+ NET019[15] WLPY_LD WLPYB_LD NET09[7] NET07[7] NET013[7] S1AHSF400W40_XDRV_LA512
XWLDV_0<8> NET05[8] NET018[8] NET017[48] NET017[49] NET017[50] NET017[51] 
+ NET017[52] NET017[53] NET04[8] NET015[56] NET015[57] NET015[58] NET015[59] 
+ NET015[60] NET015[61] NET015[62] NET011[32] NET011[33] NET011[34] NET011[35] 
+ NET012[64] NET012[65] NET012[66] NET012[67] NET012[68] NET012[69] NET012[70] 
+ NET012[71] NET014[64] NET014[65] NET014[66] NET014[67] NET014[68] NET014[69] 
+ NET014[70] NET014[71] NET03 NET016[8] NET010[8] VDDHD VDDI VSSI NET019[16] 
+ NET019[17] WLPY_LD WLPYB_LD NET09[8] NET07[8] NET013[8] S1AHSF400W40_XDRV_LA512
XWLDV_0<9> NET05[9] NET018[9] NET017[54] NET017[55] NET017[56] NET017[57] 
+ NET017[58] NET017[59] NET04[9] NET015[63] NET015[64] NET015[65] NET015[66] 
+ NET015[67] NET015[68] NET015[69] NET011[36] NET011[37] NET011[38] NET011[39] 
+ NET012[72] NET012[73] NET012[74] NET012[75] NET012[76] NET012[77] NET012[78] 
+ NET012[79] NET014[72] NET014[73] NET014[74] NET014[75] NET014[76] NET014[77] 
+ NET014[78] NET014[79] NET03 NET016[9] NET010[9] VDDHD VDDI VSSI NET019[18] 
+ NET019[19] WLPY_LD WLPYB_LD NET09[9] NET07[9] NET013[9] S1AHSF400W40_XDRV_LA512
XWLDV_0<10> NET05[10] NET018[10] NET017[60] NET017[61] NET017[62] NET017[63] 
+ NET017[64] NET017[65] NET04[10] NET015[70] NET015[71] NET015[72] NET015[73] 
+ NET015[74] NET015[75] NET015[76] NET011[40] NET011[41] NET011[42] NET011[43] 
+ NET012[80] NET012[81] NET012[82] NET012[83] NET012[84] NET012[85] NET012[86] 
+ NET012[87] NET014[80] NET014[81] NET014[82] NET014[83] NET014[84] NET014[85] 
+ NET014[86] NET014[87] NET03 NET016[10] NET010[10] VDDHD VDDI VSSI NET019[20] 
+ NET019[21] WLPY_LD WLPYB_LD NET09[10] NET07[10] NET013[10] S1AHSF400W40_XDRV_LA512
XWLDV_0<11> NET05[11] NET018[11] NET017[66] NET017[67] NET017[68] NET017[69] 
+ NET017[70] NET017[71] NET04[11] NET015[77] NET015[78] NET015[79] NET015[80] 
+ NET015[81] NET015[82] NET015[83] NET011[44] NET011[45] NET011[46] NET011[47] 
+ NET012[88] NET012[89] NET012[90] NET012[91] NET012[92] NET012[93] NET012[94] 
+ NET012[95] NET014[88] NET014[89] NET014[90] NET014[91] NET014[92] NET014[93] 
+ NET014[94] NET014[95] NET03 NET016[11] NET010[11] VDDHD VDDI VSSI NET019[22] 
+ NET019[23] WLPY_LD WLPYB_LD NET09[11] NET07[11] NET013[11] S1AHSF400W40_XDRV_LA512
XWLDV_0<12> NET05[12] NET018[12] NET017[72] NET017[73] NET017[74] NET017[75] 
+ NET017[76] NET017[77] NET04[12] NET015[84] NET015[85] NET015[86] NET015[87] 
+ NET015[88] NET015[89] NET015[90] NET011[48] NET011[49] NET011[50] NET011[51] 
+ NET012[96] NET012[97] NET012[98] NET012[99] NET012[100] NET012[101] 
+ NET012[102] NET012[103] NET014[96] NET014[97] NET014[98] NET014[99] 
+ NET014[100] NET014[101] NET014[102] NET014[103] NET03 NET016[12] NET010[12] 
+ VDDHD VDDI VSSI NET019[24] NET019[25] WLPY_LD WLPYB_LD NET09[12] NET07[12] 
+ NET013[12] S1AHSF400W40_XDRV_LA512
XWLDV_0<13> NET05[13] NET018[13] NET017[78] NET017[79] NET017[80] NET017[81] 
+ NET017[82] NET017[83] NET04[13] NET015[91] NET015[92] NET015[93] NET015[94] 
+ NET015[95] NET015[96] NET015[97] NET011[52] NET011[53] NET011[54] NET011[55] 
+ NET012[104] NET012[105] NET012[106] NET012[107] NET012[108] NET012[109] 
+ NET012[110] NET012[111] NET014[104] NET014[105] NET014[106] NET014[107] 
+ NET014[108] NET014[109] NET014[110] NET014[111] NET03 NET016[13] NET010[13] 
+ VDDHD VDDI VSSI NET019[26] NET019[27] WLPY_LD WLPYB_LD NET09[13] NET07[13] 
+ NET013[13] S1AHSF400W40_XDRV_LA512
XWLDV_0<14> NET05[14] NET018[14] NET017[84] NET017[85] NET017[86] NET017[87] 
+ NET017[88] NET017[89] NET04[14] NET015[98] NET015[99] NET015[100] 
+ NET015[101] NET015[102] NET015[103] NET015[104] NET011[56] NET011[57] 
+ NET011[58] NET011[59] NET012[112] NET012[113] NET012[114] NET012[115] 
+ NET012[116] NET012[117] NET012[118] NET012[119] NET014[112] NET014[113] 
+ NET014[114] NET014[115] NET014[116] NET014[117] NET014[118] NET014[119] 
+ NET03 NET016[14] NET010[14] VDDHD VDDI VSSI NET019[28] NET019[29] WLPY_LD 
+ WLPYB_LD NET09[14] NET07[14] NET013[14] S1AHSF400W40_XDRV_LA512
XWLDV_0<15> NET05[15] NET018[15] NET017[90] NET017[91] NET017[92] NET017[93] 
+ NET017[94] NET017[95] NET04[15] NET015[105] NET015[106] NET015[107] 
+ NET015[108] NET015[109] NET015[110] NET015[111] NET011[60] NET011[61] 
+ NET011[62] NET011[63] NET012[120] NET012[121] NET012[122] NET012[123] 
+ NET012[124] NET012[125] NET012[126] NET012[127] NET014[120] NET014[121] 
+ NET014[122] NET014[123] NET014[124] NET014[125] NET014[126] NET014[127] 
+ NET03 NET016[15] NET010[15] VDDHD VDDI VSSI NET019[30] NET019[31] WLPY_LD 
+ WLPYB_LD NET09[15] NET07[15] NET013[15] S1AHSF400W40_XDRV_LA512
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    WLPY_LD
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_WLPY_LD VDDHD VDDI VSSI WLPYB_LD WLPY_LD
*.PININFO VDDHD:B VDDI:B VSSI:B WLPYB_LD:B WLPY_LD:B
XI29 NET10[0] NET10[1] NET10[2] NET10[3] NET10[4] NET10[5] NET10[6] NET10[7] 
+ NET9[0] NET9[1] NET9[2] NET9[3] NET9[4] NET9[5] NET9[6] NET9[7] NET8 NET15 
+ VDDHD VDDI VSSI NET11[0] NET11[1] NET11[2] NET11[3] NET11[4] NET11[5] 
+ NET11[6] NET11[7] NET11[8] NET11[9] NET11[10] NET11[11] NET11[12] NET11[13] 
+ NET11[14] NET11[15] NET11[16] NET11[17] NET11[18] NET11[19] NET11[20] 
+ NET11[21] NET11[22] NET11[23] NET11[24] NET11[25] NET11[26] NET11[27] 
+ NET11[28] NET11[29] NET11[30] NET11[31] NET11[32] NET11[33] NET11[34] 
+ NET11[35] NET11[36] NET11[37] NET11[38] NET11[39] NET11[40] NET11[41] 
+ NET11[42] NET11[43] NET11[44] NET11[45] NET11[46] NET11[47] NET11[48] 
+ NET11[49] NET11[50] NET11[51] NET11[52] NET11[53] NET11[54] NET11[55] 
+ NET11[56] NET11[57] NET11[58] NET11[59] NET11[60] NET11[61] NET11[62] 
+ NET11[63] WLPY_LD WLPYB_LD S1AHSF400W40_WLDV_64X1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    WLPY_LD_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_WLPY_LD_SIM CVDDHD CVDDI VDDHD VDDI VSSI WLPYB_LD_BT WLPYB_LD_TP 
+ WLPY_LD_BT WLPY_LD_TP
*.PININFO CVDDHD:B CVDDI:B VDDHD:B VDDI:B VSSI:B WLPYB_LD_BT:B WLPYB_LD_TP:B 
*.PININFO WLPY_LD_BT:B WLPY_LD_TP:B
XI0 NET013 NET011 NET014 NET010 NET012 S1AHSF400W40_WLPY_32_LD
XWLPY_LD NET13 NET12 NET14 NET10 NET11 S1AHSF400W40_WLPY_LD
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_WLDV_D
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_WLDV_D DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] 
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] 
+ DEC_Y[7] PD_BUF RW_RE VDDHD VDDI VSSI WL[0] WL[1] WLPY WLPYB WLP_SAE 
+ WLP_SAE_TK YL[0]
*.PININFO WL[0]:O WL[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B PD_BUF:B RW_RE:B VDDHD:B VDDI:B VSSI:B WLPY:B WLPYB:B 
*.PININFO WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XWLDV_0 DEC_X0[0] DEC_X0[1] NET046[0] NET046[1] NET046[2] NET046[3] NET046[4] 
+ NET046[5] DEC_X1[0] NET044[0] NET044[1] NET044[2] NET044[3] NET044[4] 
+ NET044[5] NET044[6] NET040[0] NET040[1] NET040[2] NET040[3] NET041[0] 
+ NET041[1] NET041[2] NET041[3] NET041[4] NET041[5] NET041[6] NET041[7] 
+ NET043[0] NET043[1] NET043[2] NET043[3] NET043[4] NET043[5] NET043[6] 
+ NET043[7] PD_BUF NET29 NET039 VDDHD VDDI VSSI WL[0] WL[1] WLPY WLPYB NET038 
+ NET014 NET042 S1AHSF400W40_XDRV_LA512
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_WLDV_D_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_WLDV_D_SIM CVDDHD CVDDI DEC_X0_BT[0] DEC_X0_BT[1] DEC_X0_BT[2] 
+ DEC_X0_BT[3] DEC_X0_BT[4] DEC_X0_BT[5] DEC_X0_BT[6] DEC_X0_BT[7] 
+ DEC_X0_TP[0] DEC_X0_TP[1] DEC_X0_TP[2] DEC_X0_TP[3] DEC_X0_TP[4] 
+ DEC_X0_TP[5] DEC_X0_TP[6] DEC_X0_TP[7] DEC_X1_BT[0] DEC_X1_BT[1] 
+ DEC_X1_BT[2] DEC_X1_BT[3] DEC_X1_BT[4] DEC_X1_BT[5] DEC_X1_BT[6] 
+ DEC_X1_BT[7] DEC_X1_TP[0] DEC_X1_TP[1] DEC_X1_TP[2] DEC_X1_TP[3] 
+ DEC_X1_TP[4] DEC_X1_TP[5] DEC_X1_TP[6] DEC_X1_TP[7] DEC_X2_BT[0] 
+ DEC_X2_BT[1] DEC_X2_BT[2] DEC_X2_BT[3] DEC_X2_TP[0] DEC_X2_TP[1] 
+ DEC_X2_TP[2] DEC_X2_TP[3] DEC_X3_BT[0] DEC_X3_BT[1] DEC_X3_BT[2] 
+ DEC_X3_BT[3] DEC_X3_BT[4] DEC_X3_BT[5] DEC_X3_BT[6] DEC_X3_BT[7] 
+ DEC_X3_TP[0] DEC_X3_TP[1] DEC_X3_TP[2] DEC_X3_TP[3] DEC_X3_TP[4] 
+ DEC_X3_TP[5] DEC_X3_TP[6] DEC_X3_TP[7] DEC_Y_BT[0] DEC_Y_BT[1] DEC_Y_BT[2] 
+ DEC_Y_BT[3] DEC_Y_BT[4] DEC_Y_BT[5] DEC_Y_BT[6] DEC_Y_BT[7] DEC_Y_TP[0] 
+ DEC_Y_TP[1] DEC_Y_TP[2] DEC_Y_TP[3] DEC_Y_TP[4] DEC_Y_TP[5] DEC_Y_TP[6] 
+ DEC_Y_TP[7] PD_BUF_BT PD_BUF_TP PD_CVDDBUF_BT PD_CVDDBUF_TP RW_RE_BT 
+ RW_RE_TP VDDHD VDDI VSSI WLPYB_BT WLPYB_TP WLPY_BT WLPY_TP WLP_SAE_BT 
+ WLP_SAE_TK_BT WLP_SAE_TK_TP WLP_SAE_TP WL_LT[0] WL_LT[1] WL_RT[0] WL_RT[1] 
+ YL_BT[0] YL_TP[0]
*.PININFO DEC_X0_BT[0]:I DEC_X0_BT[1]:I DEC_X0_BT[2]:I DEC_X0_BT[3]:I 
*.PININFO DEC_X0_BT[4]:I DEC_X0_BT[5]:I DEC_X0_BT[6]:I DEC_X0_BT[7]:I 
*.PININFO DEC_X1_BT[0]:I DEC_X1_BT[1]:I DEC_X1_BT[2]:I DEC_X1_BT[3]:I 
*.PININFO DEC_X1_BT[4]:I DEC_X1_BT[5]:I DEC_X1_BT[6]:I DEC_X1_BT[7]:I 
*.PININFO PD_BUF_BT:I PD_CVDDBUF_BT:I RW_RE_TP:I DEC_X0_TP[0]:O DEC_X0_TP[1]:O 
*.PININFO DEC_X0_TP[2]:O DEC_X0_TP[3]:O DEC_X0_TP[4]:O DEC_X0_TP[5]:O 
*.PININFO DEC_X0_TP[6]:O DEC_X0_TP[7]:O DEC_X1_TP[0]:O DEC_X1_TP[1]:O 
*.PININFO DEC_X1_TP[2]:O DEC_X1_TP[3]:O DEC_X1_TP[4]:O DEC_X1_TP[5]:O 
*.PININFO DEC_X1_TP[6]:O DEC_X1_TP[7]:O PD_BUF_TP:O PD_CVDDBUF_TP:O CVDDHD:B 
*.PININFO CVDDI:B DEC_X2_BT[0]:B DEC_X2_BT[1]:B DEC_X2_BT[2]:B DEC_X2_BT[3]:B 
*.PININFO DEC_X2_TP[0]:B DEC_X2_TP[1]:B DEC_X2_TP[2]:B DEC_X2_TP[3]:B 
*.PININFO DEC_X3_BT[0]:B DEC_X3_BT[1]:B DEC_X3_BT[2]:B DEC_X3_BT[3]:B 
*.PININFO DEC_X3_BT[4]:B DEC_X3_BT[5]:B DEC_X3_BT[6]:B DEC_X3_BT[7]:B 
*.PININFO DEC_X3_TP[0]:B DEC_X3_TP[1]:B DEC_X3_TP[2]:B DEC_X3_TP[3]:B 
*.PININFO DEC_X3_TP[4]:B DEC_X3_TP[5]:B DEC_X3_TP[6]:B DEC_X3_TP[7]:B 
*.PININFO DEC_Y_BT[0]:B DEC_Y_BT[1]:B DEC_Y_BT[2]:B DEC_Y_BT[3]:B 
*.PININFO DEC_Y_BT[4]:B DEC_Y_BT[5]:B DEC_Y_BT[6]:B DEC_Y_BT[7]:B 
*.PININFO DEC_Y_TP[0]:B DEC_Y_TP[1]:B DEC_Y_TP[2]:B DEC_Y_TP[3]:B 
*.PININFO DEC_Y_TP[4]:B DEC_Y_TP[5]:B DEC_Y_TP[6]:B DEC_Y_TP[7]:B RW_RE_BT:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLPYB_BT:B WLPYB_TP:B WLPY_BT:B WLPY_TP:B 
*.PININFO WLP_SAE_BT:B WLP_SAE_TK_BT:B WLP_SAE_TK_TP:B WLP_SAE_TP:B WL_LT[0]:B 
*.PININFO WL_LT[1]:B WL_RT[0]:B WL_RT[1]:B YL_BT[0]:B YL_TP[0]:B
XI24 NET038[0] NET038[1] NET038[2] NET038[3] NET038[4] NET038[5] NET038[6] 
+ NET038[7] NET037[0] NET037[1] NET037[2] NET037[3] NET037[4] NET037[5] 
+ NET037[6] NET037[7] NET036[0] NET036[1] NET036[2] NET036[3] NET035[0] 
+ NET035[1] NET035[2] NET035[3] NET035[4] NET035[5] NET035[6] NET035[7] 
+ NET034[0] NET034[1] NET034[2] NET034[3] NET034[4] NET034[5] NET034[6] 
+ NET034[7] NET31 NET033 NET38 NET32 NET37 NET34[0] NET34[1] NET33 NET30 
+ NET032 NET031 NET03 S1AHSF400W40_BK_WLDV_D
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SIM_HB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SIM_HB AWT BIST BWEBM_LL BWEBM_LR BWEB_LL BWEB_LR CEB CEBM CLK DM_LL 
+ DM_LR D_LL D_LR FAD1[0] FAD1[1] FAD1[2] FAD1[3] FAD1[4] FAD1[5] FAD1[6] 
+ FAD1[7] FAD1[8] FAD1[9] FAD1[10] FAD2[0] FAD2[1] FAD2[2] FAD2[3] FAD2[4] 
+ FAD2[5] FAD2[6] FAD2[7] FAD2[8] FAD2[9] FAD2[10] PD PTSEL Q_LL Q_LR REDEN1 
+ REDEN2 RSTB RTSEL[0] RTSEL[1] SCLK SDIN SDOUT TM VDDI VSSI WEB WEBM 
+ WL_TK_ACT[0] WL_TK_ACT[1] WL_TK_ACT[2] WL_TK_ACT[3] WL_TK_ACT[4] 
+ WL_TK_ACT[5] WL_TK_ACT[6] WL_TK_ACT[7] WL_TK_ACT[8] WL_TK_ACT[9] 
+ WL_TK_ACT[10] WL_TK_ACT[11] WL_TK_ACT[12] WL_TK_ACT[13] WL_TK_ACT[14] 
+ WL_TK_ACT[15] WL_TK_ACT[16] WL_TK_ACT[17] WL_TK_ACT[18] WL_TK_ACT[19] 
+ WL_TK_ACT[20] WL_TK_ACT[21] WL_TK_ACT[22] WL_TK_ACT[23] WL_TK_ACT[24] 
+ WL_TK_ACT[25] WL_TK_ACT[26] WL_TK_ACT[27] WL_TK_ACT[28] WL_TK_ACT[29] 
+ WL_TK_ACT[30] WL_TK_ACT[31] WL_TK_ACT[32] WL_TK_ACT[33] WL_TK_ACT[34] 
+ WL_TK_ACT[35] WL_TK_ACT[36] WL_TK_ACT[37] WL_TK_ACT[38] WL_TK_ACT[39] 
+ WL_TK_ACT[40] WL_TK_ACT[41] WL_TK_ACT[42] WL_TK_ACT[43] WL_TK_ACT[44] 
+ WL_TK_ACT[45] WL_TK_ACT[46] WL_TK_ACT[47] WL_TK_ACT[48] WL_TK_ACT[49] 
+ WL_TK_ACT[50] WL_TK_ACT[51] WL_TK_ACT[52] WL_TK_ACT[53] WL_TK_ACT[54] 
+ WL_TK_ACT[55] WL_TK_ACT[56] WL_TK_ACT[57] WL_TK_ACT[58] WL_TK_ACT[59] 
+ WL_TK_ACT[60] WL_TK_ACT[61] WL_TK_ACT[62] WL_TK_ACT[63] WL_TK_ACT[64] 
+ WL_TK_ACT[65] WL_TK_ACT[66] WL_TK_ACT[67] WL_TK_ACT[68] WL_TK_ACT[69] 
+ WL_TK_ACT[70] WL_TK_ACT[71] WL_TK_ACT[72] WL_TK_ACT[73] WL_TK_ACT[74] 
+ WL_TK_ACT[75] WL_TK_ACT[76] WL_TK_ACT[77] WL_TK_ACT[78] WL_TK_ACT[79] 
+ WL_TK_ACT[80] WL_TK_ACT[81] WL_TK_ACT[82] WL_TK_ACT[83] WL_TK_ACT[84] 
+ WL_TK_ACT[85] WL_TK_ACT[86] WL_TK_ACT[87] WL_TK_ACT[88] WL_TK_ACT[89] 
+ WL_TK_ACT[90] WL_TK_ACT[91] WL_TK_ACT[92] WL_TK_ACT[93] WL_TK_ACT[94] 
+ WL_TK_ACT[95] WL_TK_ACT[96] WL_TK_ACT[97] WL_TK_ACT[98] WL_TK_ACT[99] 
+ WL_TK_ACT[100] WL_TK_ACT[101] WL_TK_ACT[102] WL_TK_ACT[103] WL_TK_ACT[104] 
+ WL_TK_ACT[105] WL_TK_ACT[106] WL_TK_ACT[107] WL_TK_ACT[108] WL_TK_ACT[109] 
+ WL_TK_ACT[110] WL_TK_ACT[111] WL_TK_ACT[112] WL_TK_ACT[113] WL_TK_ACT[114] 
+ WL_TK_ACT[115] WL_TK_ACT[116] WL_TK_ACT[117] WL_TK_ACT[118] WL_TK_ACT[119] 
+ WL_TK_ACT[120] WL_TK_ACT[121] WL_TK_ACT[122] WL_TK_ACT[123] WL_TK_ACT[124] 
+ WL_TK_ACT[125] WL_TK_ACT[126] WL_TK_ACT[127] WL_TK_ACT[128] WL_TK_ACT[129] 
+ WL_TK_ACT[130] WL_TK_ACT[131] WL_TK_ACT[132] WL_TK_ACT[133] WL_TK_ACT[134] 
+ WL_TK_ACT[135] WL_TK_ACT[136] WL_TK_ACT[137] WL_TK_ACT[138] WL_TK_ACT[139] 
+ WL_TK_ACT[140] WL_TK_ACT[141] WL_TK_ACT[142] WL_TK_ACT[143] WL_TK_ACT[144] 
+ WL_TK_ACT[145] WL_TK_ACT[146] WL_TK_ACT[147] WL_TK_ACT[148] WL_TK_ACT[149] 
+ WL_TK_ACT[150] WL_TK_ACT[151] WL_TK_ACT[152] WL_TK_ACT[153] WL_TK_ACT[154] 
+ WL_TK_ACT[155] WL_TK_ACT[156] WL_TK_ACT[157] WL_TK_ACT[158] WL_TK_ACT[159] 
+ WL_TK_ACT[160] WL_TK_ACT[161] WL_TK_ACT[162] WL_TK_ACT[163] WL_TK_ACT[164] 
+ WL_TK_ACT[165] WL_TK_ACT[166] WL_TK_ACT[167] WL_TK_ACT[168] WL_TK_ACT[169] 
+ WL_TK_ACT[170] WL_TK_ACT[171] WL_TK_ACT[172] WL_TK_ACT[173] WL_TK_ACT[174] 
+ WL_TK_ACT[175] WL_TK_ACT[176] WL_TK_ACT[177] WL_TK_ACT[178] WL_TK_ACT[179] 
+ WL_TK_ACT[180] WL_TK_ACT[181] WL_TK_ACT[182] WL_TK_ACT[183] WL_TK_ACT[184] 
+ WL_TK_ACT[185] WL_TK_ACT[186] WL_TK_ACT[187] WL_TK_ACT[188] WL_TK_ACT[189] 
+ WL_TK_ACT[190] WL_TK_ACT[191] WL_TK_ACT[192] WL_TK_ACT[193] WL_TK_ACT[194] 
+ WL_TK_ACT[195] WL_TK_ACT[196] WL_TK_ACT[197] WL_TK_ACT[198] WL_TK_ACT[199] 
+ WL_TK_ACT[200] WL_TK_ACT[201] WL_TK_ACT[202] WL_TK_ACT[203] WL_TK_ACT[204] 
+ WL_TK_ACT[205] WL_TK_ACT[206] WL_TK_ACT[207] WL_TK_ACT[208] WL_TK_ACT[209] 
+ WL_TK_ACT[210] WL_TK_ACT[211] WL_TK_ACT[212] WL_TK_ACT[213] WL_TK_ACT[214] 
+ WL_TK_ACT[215] WL_TK_ACT[216] WL_TK_ACT[217] WL_TK_ACT[218] WL_TK_ACT[219] 
+ WL_TK_ACT[220] WL_TK_ACT[221] WL_TK_ACT[222] WL_TK_ACT[223] WL_TK_ACT[224] 
+ WL_TK_ACT[225] WL_TK_ACT[226] WL_TK_ACT[227] WL_TK_ACT[228] WL_TK_ACT[229] 
+ WL_TK_ACT[230] WL_TK_ACT[231] WL_TK_ACT[232] WL_TK_ACT[233] WL_TK_ACT[234] 
+ WL_TK_ACT[235] WL_TK_ACT[236] WL_TK_ACT[237] WL_TK_ACT[238] WL_TK_ACT[239] 
+ WL_TK_ACT[240] WL_TK_ACT[241] WL_TK_ACT[242] WL_TK_ACT[243] WL_TK_ACT[244] 
+ WL_TK_ACT[245] WL_TK_ACT[246] WL_TK_ACT[247] WL_TK_ACT[248] WL_TK_ACT[249] 
+ WL_TK_ACT[250] WL_TK_ACT[251] WL_TK_ACT[252] WL_TK_ACT[253] WL_TK_ACT[254] 
+ WL_TK_ACT[255] WL_TK_ACT[256] WL_TK_ACT[257] WL_TK_ACT[258] WL_TK_ACT[259] 
+ WL_TK_ACT[260] WL_TK_ACT[261] WL_TK_ACT[262] WL_TK_ACT[263] WL_TK_ACT[264] 
+ WL_TK_ACT[265] WL_TK_ACT[266] WL_TK_ACT[267] WL_TK_ACT[268] WL_TK_ACT[269] 
+ WL_TK_ACT[270] WL_TK_ACT[271] WL_TK_ACT[272] WL_TK_ACT[273] WL_TK_ACT[274] 
+ WL_TK_ACT[275] WL_TK_ACT[276] WL_TK_ACT[277] WL_TK_ACT[278] WL_TK_ACT[279] 
+ WL_TK_ACT[280] WL_TK_ACT[281] WL_TK_ACT[282] WL_TK_ACT[283] WL_TK_ACT[284] 
+ WL_TK_ACT[285] WL_TK_ACT[286] WL_TK_ACT[287] WL_TK_ACT[288] WL_TK_ACT[289] 
+ WL_TK_ACT[290] WL_TK_ACT[291] WL_TK_ACT[292] WL_TK_ACT[293] WL_TK_ACT[294] 
+ WL_TK_ACT[295] WL_TK_ACT[296] WL_TK_ACT[297] WL_TK_ACT[298] WL_TK_ACT[299] 
+ WL_TK_ACT[300] WL_TK_ACT[301] WL_TK_ACT[302] WL_TK_ACT[303] WL_TK_ACT[304] 
+ WL_TK_ACT[305] WL_TK_ACT[306] WL_TK_ACT[307] WL_TK_ACT[308] WL_TK_ACT[309] 
+ WL_TK_ACT[310] WL_TK_ACT[311] WL_TK_ACT[312] WL_TK_ACT[313] WL_TK_ACT[314] 
+ WL_TK_ACT[315] WL_TK_ACT[316] WL_TK_ACT[317] WL_TK_ACT[318] WL_TK_ACT[319] 
+ WL_TK_ACT[320] WL_TK_ACT[321] WL_TK_ACT[322] WL_TK_ACT[323] WL_TK_ACT[324] 
+ WL_TK_ACT[325] WL_TK_ACT[326] WL_TK_ACT[327] WL_TK_ACT[328] WL_TK_ACT[329] 
+ WL_TK_ACT[330] WL_TK_ACT[331] WL_TK_ACT[332] WL_TK_ACT[333] WL_TK_ACT[334] 
+ WL_TK_ACT[335] WL_TK_ACT[336] WL_TK_ACT[337] WL_TK_ACT[338] WL_TK_ACT[339] 
+ WL_TK_ACT[340] WL_TK_ACT[341] WL_TK_ACT[342] WL_TK_ACT[343] WL_TK_ACT[344] 
+ WL_TK_ACT[345] WL_TK_ACT[346] WL_TK_ACT[347] WL_TK_ACT[348] WL_TK_ACT[349] 
+ WL_TK_ACT[350] WL_TK_ACT[351] WL_TK_ACT[352] WL_TK_ACT[353] WL_TK_ACT[354] 
+ WL_TK_ACT[355] WL_TK_ACT[356] WL_TK_ACT[357] WL_TK_ACT[358] WL_TK_ACT[359] 
+ WL_TK_ACT[360] WL_TK_ACT[361] WL_TK_ACT[362] WL_TK_ACT[363] WL_TK_ACT[364] 
+ WL_TK_ACT[365] WL_TK_ACT[366] WL_TK_ACT[367] WL_TK_ACT[368] WL_TK_ACT[369] 
+ WL_TK_ACT[370] WL_TK_ACT[371] WL_TK_ACT[372] WL_TK_ACT[373] WL_TK_ACT[374] 
+ WL_TK_ACT[375] WL_TK_ACT[376] WL_TK_ACT[377] WL_TK_ACT[378] WL_TK_ACT[379] 
+ WL_TK_ACT[380] WL_TK_ACT[381] WL_TK_ACT[382] WL_TK_ACT[383] WL_TK_ACT[384] 
+ WL_TK_ACT[385] WL_TK_ACT[386] WL_TK_ACT[387] WL_TK_ACT[388] WL_TK_ACT[389] 
+ WL_TK_ACT[390] WL_TK_ACT[391] WL_TK_ACT[392] WL_TK_ACT[393] WL_TK_ACT[394] 
+ WL_TK_ACT[395] WL_TK_ACT[396] WL_TK_ACT[397] WL_TK_ACT[398] WL_TK_ACT[399] 
+ WL_TK_ACT[400] WL_TK_ACT[401] WL_TK_ACT[402] WL_TK_ACT[403] WL_TK_ACT[404] 
+ WL_TK_ACT[405] WL_TK_ACT[406] WL_TK_ACT[407] WL_TK_ACT[408] WL_TK_ACT[409] 
+ WL_TK_ACT[410] WL_TK_ACT[411] WL_TK_ACT[412] WL_TK_ACT[413] WL_TK_ACT[414] 
+ WL_TK_ACT[415] WL_TK_ACT[416] WL_TK_ACT[417] WL_TK_ACT[418] WL_TK_ACT[419] 
+ WL_TK_ACT[420] WL_TK_ACT[421] WL_TK_ACT[422] WL_TK_ACT[423] WL_TK_ACT[424] 
+ WL_TK_ACT[425] WL_TK_ACT[426] WL_TK_ACT[427] WL_TK_ACT[428] WL_TK_ACT[429] 
+ WL_TK_ACT[430] WL_TK_ACT[431] WL_TK_ACT[432] WL_TK_ACT[433] WL_TK_ACT[434] 
+ WL_TK_ACT[435] WL_TK_ACT[436] WL_TK_ACT[437] WL_TK_ACT[438] WL_TK_ACT[439] 
+ WL_TK_ACT[440] WL_TK_ACT[441] WL_TK_ACT[442] WL_TK_ACT[443] WL_TK_ACT[444] 
+ WL_TK_ACT[445] WL_TK_ACT[446] WL_TK_ACT[447] WL_TK_ACT[448] WL_TK_ACT[449] 
+ WL_TK_ACT[450] WL_TK_ACT[451] WL_TK_ACT[452] WL_TK_ACT[453] WL_TK_ACT[454] 
+ WL_TK_ACT[455] WL_TK_ACT[456] WL_TK_ACT[457] WL_TK_ACT[458] WL_TK_ACT[459] 
+ WL_TK_ACT[460] WL_TK_ACT[461] WL_TK_ACT[462] WL_TK_ACT[463] WL_TK_ACT[464] 
+ WL_TK_ACT[465] WL_TK_ACT[466] WL_TK_ACT[467] WL_TK_ACT[468] WL_TK_ACT[469] 
+ WL_TK_ACT[470] WL_TK_ACT[471] WL_TK_ACT[472] WL_TK_ACT[473] WL_TK_ACT[474] 
+ WL_TK_ACT[475] WL_TK_ACT[476] WL_TK_ACT[477] WL_TK_ACT[478] WL_TK_ACT[479] 
+ WL_TK_ACT[480] WL_TK_ACT[481] WL_TK_ACT[482] WL_TK_ACT[483] WL_TK_ACT[484] 
+ WL_TK_ACT[485] WL_TK_ACT[486] WL_TK_ACT[487] WL_TK_ACT[488] WL_TK_ACT[489] 
+ WL_TK_ACT[490] WL_TK_ACT[491] WL_TK_ACT[492] WL_TK_ACT[493] WL_TK_ACT[494] 
+ WL_TK_ACT[495] WL_TK_ACT[496] WL_TK_ACT[497] WL_TK_ACT[498] WL_TK_ACT[499] 
+ WL_TK_ACT[500] WL_TK_ACT[501] WL_TK_ACT[502] WL_TK_ACT[503] WL_TK_ACT[504] 
+ WL_TK_ACT[505] WL_TK_ACT[506] WL_TK_ACT[507] WL_TK_ACT[508] WL_TK_ACT[509] 
+ WL_TK_ACT[510] WL_TK_ACT[511] WL_TK_LD WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] 
+ X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] 
+ XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YM[0] YM[1] YM[2] 
+ YM[3]
*.PININFO AWT:I BIST:I BWEBM_LL:I BWEBM_LR:I BWEB_LL:I BWEB_LR:I CEB:I CEBM:I 
*.PININFO CLK:I DM_LL:I DM_LR:I D_LL:I D_LR:I FAD1[0]:I FAD1[1]:I FAD1[2]:I 
*.PININFO FAD1[3]:I FAD1[4]:I FAD1[5]:I FAD1[6]:I FAD1[7]:I FAD1[8]:I 
*.PININFO FAD1[9]:I FAD1[10]:I FAD2[0]:I FAD2[1]:I FAD2[2]:I FAD2[3]:I 
*.PININFO FAD2[4]:I FAD2[5]:I FAD2[6]:I FAD2[7]:I FAD2[8]:I FAD2[9]:I 
*.PININFO FAD2[10]:I PD:I PTSEL:I REDEN1:I REDEN2:I RSTB:I RTSEL[0]:I 
*.PININFO RTSEL[1]:I SCLK:I SDIN:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I 
*.PININFO XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I 
*.PININFO Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I Q_LL:O Q_LR:O SDOUT:O 
*.PININFO VDDI:B VSSI:B WL_TK_ACT[0]:B WL_TK_ACT[1]:B WL_TK_ACT[2]:B 
*.PININFO WL_TK_ACT[3]:B WL_TK_ACT[4]:B WL_TK_ACT[5]:B WL_TK_ACT[6]:B 
*.PININFO WL_TK_ACT[7]:B WL_TK_ACT[8]:B WL_TK_ACT[9]:B WL_TK_ACT[10]:B 
*.PININFO WL_TK_ACT[11]:B WL_TK_ACT[12]:B WL_TK_ACT[13]:B WL_TK_ACT[14]:B 
*.PININFO WL_TK_ACT[15]:B WL_TK_ACT[16]:B WL_TK_ACT[17]:B WL_TK_ACT[18]:B 
*.PININFO WL_TK_ACT[19]:B WL_TK_ACT[20]:B WL_TK_ACT[21]:B WL_TK_ACT[22]:B 
*.PININFO WL_TK_ACT[23]:B WL_TK_ACT[24]:B WL_TK_ACT[25]:B WL_TK_ACT[26]:B 
*.PININFO WL_TK_ACT[27]:B WL_TK_ACT[28]:B WL_TK_ACT[29]:B WL_TK_ACT[30]:B 
*.PININFO WL_TK_ACT[31]:B WL_TK_ACT[32]:B WL_TK_ACT[33]:B WL_TK_ACT[34]:B 
*.PININFO WL_TK_ACT[35]:B WL_TK_ACT[36]:B WL_TK_ACT[37]:B WL_TK_ACT[38]:B 
*.PININFO WL_TK_ACT[39]:B WL_TK_ACT[40]:B WL_TK_ACT[41]:B WL_TK_ACT[42]:B 
*.PININFO WL_TK_ACT[43]:B WL_TK_ACT[44]:B WL_TK_ACT[45]:B WL_TK_ACT[46]:B 
*.PININFO WL_TK_ACT[47]:B WL_TK_ACT[48]:B WL_TK_ACT[49]:B WL_TK_ACT[50]:B 
*.PININFO WL_TK_ACT[51]:B WL_TK_ACT[52]:B WL_TK_ACT[53]:B WL_TK_ACT[54]:B 
*.PININFO WL_TK_ACT[55]:B WL_TK_ACT[56]:B WL_TK_ACT[57]:B WL_TK_ACT[58]:B 
*.PININFO WL_TK_ACT[59]:B WL_TK_ACT[60]:B WL_TK_ACT[61]:B WL_TK_ACT[62]:B 
*.PININFO WL_TK_ACT[63]:B WL_TK_ACT[64]:B WL_TK_ACT[65]:B WL_TK_ACT[66]:B 
*.PININFO WL_TK_ACT[67]:B WL_TK_ACT[68]:B WL_TK_ACT[69]:B WL_TK_ACT[70]:B 
*.PININFO WL_TK_ACT[71]:B WL_TK_ACT[72]:B WL_TK_ACT[73]:B WL_TK_ACT[74]:B 
*.PININFO WL_TK_ACT[75]:B WL_TK_ACT[76]:B WL_TK_ACT[77]:B WL_TK_ACT[78]:B 
*.PININFO WL_TK_ACT[79]:B WL_TK_ACT[80]:B WL_TK_ACT[81]:B WL_TK_ACT[82]:B 
*.PININFO WL_TK_ACT[83]:B WL_TK_ACT[84]:B WL_TK_ACT[85]:B WL_TK_ACT[86]:B 
*.PININFO WL_TK_ACT[87]:B WL_TK_ACT[88]:B WL_TK_ACT[89]:B WL_TK_ACT[90]:B 
*.PININFO WL_TK_ACT[91]:B WL_TK_ACT[92]:B WL_TK_ACT[93]:B WL_TK_ACT[94]:B 
*.PININFO WL_TK_ACT[95]:B WL_TK_ACT[96]:B WL_TK_ACT[97]:B WL_TK_ACT[98]:B 
*.PININFO WL_TK_ACT[99]:B WL_TK_ACT[100]:B WL_TK_ACT[101]:B WL_TK_ACT[102]:B 
*.PININFO WL_TK_ACT[103]:B WL_TK_ACT[104]:B WL_TK_ACT[105]:B WL_TK_ACT[106]:B 
*.PININFO WL_TK_ACT[107]:B WL_TK_ACT[108]:B WL_TK_ACT[109]:B WL_TK_ACT[110]:B 
*.PININFO WL_TK_ACT[111]:B WL_TK_ACT[112]:B WL_TK_ACT[113]:B WL_TK_ACT[114]:B 
*.PININFO WL_TK_ACT[115]:B WL_TK_ACT[116]:B WL_TK_ACT[117]:B WL_TK_ACT[118]:B 
*.PININFO WL_TK_ACT[119]:B WL_TK_ACT[120]:B WL_TK_ACT[121]:B WL_TK_ACT[122]:B 
*.PININFO WL_TK_ACT[123]:B WL_TK_ACT[124]:B WL_TK_ACT[125]:B WL_TK_ACT[126]:B 
*.PININFO WL_TK_ACT[127]:B WL_TK_ACT[128]:B WL_TK_ACT[129]:B WL_TK_ACT[130]:B 
*.PININFO WL_TK_ACT[131]:B WL_TK_ACT[132]:B WL_TK_ACT[133]:B WL_TK_ACT[134]:B 
*.PININFO WL_TK_ACT[135]:B WL_TK_ACT[136]:B WL_TK_ACT[137]:B WL_TK_ACT[138]:B 
*.PININFO WL_TK_ACT[139]:B WL_TK_ACT[140]:B WL_TK_ACT[141]:B WL_TK_ACT[142]:B 
*.PININFO WL_TK_ACT[143]:B WL_TK_ACT[144]:B WL_TK_ACT[145]:B WL_TK_ACT[146]:B 
*.PININFO WL_TK_ACT[147]:B WL_TK_ACT[148]:B WL_TK_ACT[149]:B WL_TK_ACT[150]:B 
*.PININFO WL_TK_ACT[151]:B WL_TK_ACT[152]:B WL_TK_ACT[153]:B WL_TK_ACT[154]:B 
*.PININFO WL_TK_ACT[155]:B WL_TK_ACT[156]:B WL_TK_ACT[157]:B WL_TK_ACT[158]:B 
*.PININFO WL_TK_ACT[159]:B WL_TK_ACT[160]:B WL_TK_ACT[161]:B WL_TK_ACT[162]:B 
*.PININFO WL_TK_ACT[163]:B WL_TK_ACT[164]:B WL_TK_ACT[165]:B WL_TK_ACT[166]:B 
*.PININFO WL_TK_ACT[167]:B WL_TK_ACT[168]:B WL_TK_ACT[169]:B WL_TK_ACT[170]:B 
*.PININFO WL_TK_ACT[171]:B WL_TK_ACT[172]:B WL_TK_ACT[173]:B WL_TK_ACT[174]:B 
*.PININFO WL_TK_ACT[175]:B WL_TK_ACT[176]:B WL_TK_ACT[177]:B WL_TK_ACT[178]:B 
*.PININFO WL_TK_ACT[179]:B WL_TK_ACT[180]:B WL_TK_ACT[181]:B WL_TK_ACT[182]:B 
*.PININFO WL_TK_ACT[183]:B WL_TK_ACT[184]:B WL_TK_ACT[185]:B WL_TK_ACT[186]:B 
*.PININFO WL_TK_ACT[187]:B WL_TK_ACT[188]:B WL_TK_ACT[189]:B WL_TK_ACT[190]:B 
*.PININFO WL_TK_ACT[191]:B WL_TK_ACT[192]:B WL_TK_ACT[193]:B WL_TK_ACT[194]:B 
*.PININFO WL_TK_ACT[195]:B WL_TK_ACT[196]:B WL_TK_ACT[197]:B WL_TK_ACT[198]:B 
*.PININFO WL_TK_ACT[199]:B WL_TK_ACT[200]:B WL_TK_ACT[201]:B WL_TK_ACT[202]:B 
*.PININFO WL_TK_ACT[203]:B WL_TK_ACT[204]:B WL_TK_ACT[205]:B WL_TK_ACT[206]:B 
*.PININFO WL_TK_ACT[207]:B WL_TK_ACT[208]:B WL_TK_ACT[209]:B WL_TK_ACT[210]:B 
*.PININFO WL_TK_ACT[211]:B WL_TK_ACT[212]:B WL_TK_ACT[213]:B WL_TK_ACT[214]:B 
*.PININFO WL_TK_ACT[215]:B WL_TK_ACT[216]:B WL_TK_ACT[217]:B WL_TK_ACT[218]:B 
*.PININFO WL_TK_ACT[219]:B WL_TK_ACT[220]:B WL_TK_ACT[221]:B WL_TK_ACT[222]:B 
*.PININFO WL_TK_ACT[223]:B WL_TK_ACT[224]:B WL_TK_ACT[225]:B WL_TK_ACT[226]:B 
*.PININFO WL_TK_ACT[227]:B WL_TK_ACT[228]:B WL_TK_ACT[229]:B WL_TK_ACT[230]:B 
*.PININFO WL_TK_ACT[231]:B WL_TK_ACT[232]:B WL_TK_ACT[233]:B WL_TK_ACT[234]:B 
*.PININFO WL_TK_ACT[235]:B WL_TK_ACT[236]:B WL_TK_ACT[237]:B WL_TK_ACT[238]:B 
*.PININFO WL_TK_ACT[239]:B WL_TK_ACT[240]:B WL_TK_ACT[241]:B WL_TK_ACT[242]:B 
*.PININFO WL_TK_ACT[243]:B WL_TK_ACT[244]:B WL_TK_ACT[245]:B WL_TK_ACT[246]:B 
*.PININFO WL_TK_ACT[247]:B WL_TK_ACT[248]:B WL_TK_ACT[249]:B WL_TK_ACT[250]:B 
*.PININFO WL_TK_ACT[251]:B WL_TK_ACT[252]:B WL_TK_ACT[253]:B WL_TK_ACT[254]:B 
*.PININFO WL_TK_ACT[255]:B WL_TK_ACT[256]:B WL_TK_ACT[257]:B WL_TK_ACT[258]:B 
*.PININFO WL_TK_ACT[259]:B WL_TK_ACT[260]:B WL_TK_ACT[261]:B WL_TK_ACT[262]:B 
*.PININFO WL_TK_ACT[263]:B WL_TK_ACT[264]:B WL_TK_ACT[265]:B WL_TK_ACT[266]:B 
*.PININFO WL_TK_ACT[267]:B WL_TK_ACT[268]:B WL_TK_ACT[269]:B WL_TK_ACT[270]:B 
*.PININFO WL_TK_ACT[271]:B WL_TK_ACT[272]:B WL_TK_ACT[273]:B WL_TK_ACT[274]:B 
*.PININFO WL_TK_ACT[275]:B WL_TK_ACT[276]:B WL_TK_ACT[277]:B WL_TK_ACT[278]:B 
*.PININFO WL_TK_ACT[279]:B WL_TK_ACT[280]:B WL_TK_ACT[281]:B WL_TK_ACT[282]:B 
*.PININFO WL_TK_ACT[283]:B WL_TK_ACT[284]:B WL_TK_ACT[285]:B WL_TK_ACT[286]:B 
*.PININFO WL_TK_ACT[287]:B WL_TK_ACT[288]:B WL_TK_ACT[289]:B WL_TK_ACT[290]:B 
*.PININFO WL_TK_ACT[291]:B WL_TK_ACT[292]:B WL_TK_ACT[293]:B WL_TK_ACT[294]:B 
*.PININFO WL_TK_ACT[295]:B WL_TK_ACT[296]:B WL_TK_ACT[297]:B WL_TK_ACT[298]:B 
*.PININFO WL_TK_ACT[299]:B WL_TK_ACT[300]:B WL_TK_ACT[301]:B WL_TK_ACT[302]:B 
*.PININFO WL_TK_ACT[303]:B WL_TK_ACT[304]:B WL_TK_ACT[305]:B WL_TK_ACT[306]:B 
*.PININFO WL_TK_ACT[307]:B WL_TK_ACT[308]:B WL_TK_ACT[309]:B WL_TK_ACT[310]:B 
*.PININFO WL_TK_ACT[311]:B WL_TK_ACT[312]:B WL_TK_ACT[313]:B WL_TK_ACT[314]:B 
*.PININFO WL_TK_ACT[315]:B WL_TK_ACT[316]:B WL_TK_ACT[317]:B WL_TK_ACT[318]:B 
*.PININFO WL_TK_ACT[319]:B WL_TK_ACT[320]:B WL_TK_ACT[321]:B WL_TK_ACT[322]:B 
*.PININFO WL_TK_ACT[323]:B WL_TK_ACT[324]:B WL_TK_ACT[325]:B WL_TK_ACT[326]:B 
*.PININFO WL_TK_ACT[327]:B WL_TK_ACT[328]:B WL_TK_ACT[329]:B WL_TK_ACT[330]:B 
*.PININFO WL_TK_ACT[331]:B WL_TK_ACT[332]:B WL_TK_ACT[333]:B WL_TK_ACT[334]:B 
*.PININFO WL_TK_ACT[335]:B WL_TK_ACT[336]:B WL_TK_ACT[337]:B WL_TK_ACT[338]:B 
*.PININFO WL_TK_ACT[339]:B WL_TK_ACT[340]:B WL_TK_ACT[341]:B WL_TK_ACT[342]:B 
*.PININFO WL_TK_ACT[343]:B WL_TK_ACT[344]:B WL_TK_ACT[345]:B WL_TK_ACT[346]:B 
*.PININFO WL_TK_ACT[347]:B WL_TK_ACT[348]:B WL_TK_ACT[349]:B WL_TK_ACT[350]:B 
*.PININFO WL_TK_ACT[351]:B WL_TK_ACT[352]:B WL_TK_ACT[353]:B WL_TK_ACT[354]:B 
*.PININFO WL_TK_ACT[355]:B WL_TK_ACT[356]:B WL_TK_ACT[357]:B WL_TK_ACT[358]:B 
*.PININFO WL_TK_ACT[359]:B WL_TK_ACT[360]:B WL_TK_ACT[361]:B WL_TK_ACT[362]:B 
*.PININFO WL_TK_ACT[363]:B WL_TK_ACT[364]:B WL_TK_ACT[365]:B WL_TK_ACT[366]:B 
*.PININFO WL_TK_ACT[367]:B WL_TK_ACT[368]:B WL_TK_ACT[369]:B WL_TK_ACT[370]:B 
*.PININFO WL_TK_ACT[371]:B WL_TK_ACT[372]:B WL_TK_ACT[373]:B WL_TK_ACT[374]:B 
*.PININFO WL_TK_ACT[375]:B WL_TK_ACT[376]:B WL_TK_ACT[377]:B WL_TK_ACT[378]:B 
*.PININFO WL_TK_ACT[379]:B WL_TK_ACT[380]:B WL_TK_ACT[381]:B WL_TK_ACT[382]:B 
*.PININFO WL_TK_ACT[383]:B WL_TK_ACT[384]:B WL_TK_ACT[385]:B WL_TK_ACT[386]:B 
*.PININFO WL_TK_ACT[387]:B WL_TK_ACT[388]:B WL_TK_ACT[389]:B WL_TK_ACT[390]:B 
*.PININFO WL_TK_ACT[391]:B WL_TK_ACT[392]:B WL_TK_ACT[393]:B WL_TK_ACT[394]:B 
*.PININFO WL_TK_ACT[395]:B WL_TK_ACT[396]:B WL_TK_ACT[397]:B WL_TK_ACT[398]:B 
*.PININFO WL_TK_ACT[399]:B WL_TK_ACT[400]:B WL_TK_ACT[401]:B WL_TK_ACT[402]:B 
*.PININFO WL_TK_ACT[403]:B WL_TK_ACT[404]:B WL_TK_ACT[405]:B WL_TK_ACT[406]:B 
*.PININFO WL_TK_ACT[407]:B WL_TK_ACT[408]:B WL_TK_ACT[409]:B WL_TK_ACT[410]:B 
*.PININFO WL_TK_ACT[411]:B WL_TK_ACT[412]:B WL_TK_ACT[413]:B WL_TK_ACT[414]:B 
*.PININFO WL_TK_ACT[415]:B WL_TK_ACT[416]:B WL_TK_ACT[417]:B WL_TK_ACT[418]:B 
*.PININFO WL_TK_ACT[419]:B WL_TK_ACT[420]:B WL_TK_ACT[421]:B WL_TK_ACT[422]:B 
*.PININFO WL_TK_ACT[423]:B WL_TK_ACT[424]:B WL_TK_ACT[425]:B WL_TK_ACT[426]:B 
*.PININFO WL_TK_ACT[427]:B WL_TK_ACT[428]:B WL_TK_ACT[429]:B WL_TK_ACT[430]:B 
*.PININFO WL_TK_ACT[431]:B WL_TK_ACT[432]:B WL_TK_ACT[433]:B WL_TK_ACT[434]:B 
*.PININFO WL_TK_ACT[435]:B WL_TK_ACT[436]:B WL_TK_ACT[437]:B WL_TK_ACT[438]:B 
*.PININFO WL_TK_ACT[439]:B WL_TK_ACT[440]:B WL_TK_ACT[441]:B WL_TK_ACT[442]:B 
*.PININFO WL_TK_ACT[443]:B WL_TK_ACT[444]:B WL_TK_ACT[445]:B WL_TK_ACT[446]:B 
*.PININFO WL_TK_ACT[447]:B WL_TK_ACT[448]:B WL_TK_ACT[449]:B WL_TK_ACT[450]:B 
*.PININFO WL_TK_ACT[451]:B WL_TK_ACT[452]:B WL_TK_ACT[453]:B WL_TK_ACT[454]:B 
*.PININFO WL_TK_ACT[455]:B WL_TK_ACT[456]:B WL_TK_ACT[457]:B WL_TK_ACT[458]:B 
*.PININFO WL_TK_ACT[459]:B WL_TK_ACT[460]:B WL_TK_ACT[461]:B WL_TK_ACT[462]:B 
*.PININFO WL_TK_ACT[463]:B WL_TK_ACT[464]:B WL_TK_ACT[465]:B WL_TK_ACT[466]:B 
*.PININFO WL_TK_ACT[467]:B WL_TK_ACT[468]:B WL_TK_ACT[469]:B WL_TK_ACT[470]:B 
*.PININFO WL_TK_ACT[471]:B WL_TK_ACT[472]:B WL_TK_ACT[473]:B WL_TK_ACT[474]:B 
*.PININFO WL_TK_ACT[475]:B WL_TK_ACT[476]:B WL_TK_ACT[477]:B WL_TK_ACT[478]:B 
*.PININFO WL_TK_ACT[479]:B WL_TK_ACT[480]:B WL_TK_ACT[481]:B WL_TK_ACT[482]:B 
*.PININFO WL_TK_ACT[483]:B WL_TK_ACT[484]:B WL_TK_ACT[485]:B WL_TK_ACT[486]:B 
*.PININFO WL_TK_ACT[487]:B WL_TK_ACT[488]:B WL_TK_ACT[489]:B WL_TK_ACT[490]:B 
*.PININFO WL_TK_ACT[491]:B WL_TK_ACT[492]:B WL_TK_ACT[493]:B WL_TK_ACT[494]:B 
*.PININFO WL_TK_ACT[495]:B WL_TK_ACT[496]:B WL_TK_ACT[497]:B WL_TK_ACT[498]:B 
*.PININFO WL_TK_ACT[499]:B WL_TK_ACT[500]:B WL_TK_ACT[501]:B WL_TK_ACT[502]:B 
*.PININFO WL_TK_ACT[503]:B WL_TK_ACT[504]:B WL_TK_ACT[505]:B WL_TK_ACT[506]:B 
*.PININFO WL_TK_ACT[507]:B WL_TK_ACT[508]:B WL_TK_ACT[509]:B WL_TK_ACT[510]:B 
*.PININFO WL_TK_ACT[511]:B WL_TK_LD:B
XCNT AWT AWT2_L1 BIST BIST2IO_L1 WL_TK CEB CEBM CKD_L1 CLK VDDHD VDDI 
+ DEC_X0_1[0] DEC_X0_1[1] DEC_X0_1[2] DEC_X0_1[3] DEC_X0_1[4] DEC_X0_1[5] 
+ DEC_X0_1[6] DEC_X0_1[7] DEC_X1_1[0] DEC_X1_1[1] DEC_X1_1[2] DEC_X1_1[3] 
+ DEC_X1_1[4] DEC_X1_1[5] DEC_X1_1[6] DEC_X1_1[7] DEC_X2_1[0] DEC_X2_1[1] 
+ DEC_X2_1[2] DEC_X2_1[3] DEC_X3_1[0] DEC_X3_1[1] DEC_X3_1[2] DEC_X3_1[3] 
+ DEC_X3_1[4] DEC_X3_1[5] DEC_X3_1[6] DEC_X3_1[7] DEC_Y_1[0] DEC_Y_1[1] 
+ DEC_Y_1[2] DEC_Y_1[3] DEC_Y_1[4] DEC_Y_1[5] DEC_Y_1[6] DEC_Y_1[7] FAD1[0] 
+ FAD1[1] FAD1[2] FAD1[3] FAD1[4] FAD1[5] FAD1[6] FAD1[7] FAD1[8] FAD1[9] 
+ FAD1[10] FAD2[0] FAD2[1] FAD2[2] FAD2[3] FAD2[4] FAD2[5] FAD2[6] FAD2[7] 
+ FAD2[8] FAD2[9] FAD2[10] NET154[0] NET154[1] PD PD_BUF_1 PD_CVDDBUF_1 PTSEL 
+ REDEN_BT REDEN1 REDEN2 REDENB_BT RSTB RTSEL[0] RTSEL[1] RW_RE_1 SCLK SDIN 
+ SDOUT TK TM TRKBL VDDHD VDDI VHI_LT VLO_LT VSSI WEB WEBM WLP_SAE_1 
+ WLP_SAEB_L1 WLP_SAE_TK_1 WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] 
+ X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] 
+ XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL_1[0] YM[0] YM[1] YM[2] YM[3] 
+ S1AHSF400W40_CNT_SIM
XIO_LD_L AWT2_L3 AWT2_L2 BIST2IO_L3 BIST2IO_L2 CKD_L3 CKD_L2 PD_BUF_L3 
+ PD_BUF_L2 VDDHD VDDI VSSI WLP_SAEB_L3 WLP_SAEB_L2 S1AHSF400W40_IO_LD_SIM
XIO_LD_R AWT2_R2 AWT2_R3 BIST2IO_R2 BIST2IO_R3 CKD_R2 CKD_R3 PD_BUF_R2 
+ PD_BUF_R3 VDDHD VDDI VSSI WLP_SAEB_R2 WLP_SAEB_R3 S1AHSF400W40_IO_LD_SIM
XIO_LL AWT2_L4 AWT2_L3 BIST2IO_L4 BIST2IO_L3 BWEBM_LL BWEB_LL CKD_L4 CKD_L3 
+ DM_LL D_LL GBLB_LL_12 GBL_LL_12 GWB_LL_12 GW_LL_12 PD_BUF_L4 PD_BUF_L3 Q_LL 
+ VDDHD VDDI VSSI WLP_SAEB_L4 WLP_SAEB_L3 S1AHSF400W40_IO_SIM
XIO_RL AWT2_L1 AWT2_R2 BIST2IO_L1 BIST2IO_R2 NET231 NET232 CKD_L1 CKD_R2 
+ NET229 NET228 NET392 NET235 NET233 NET234 PD_BUF_1 PD_BUF_R2 NET227 VDDHD 
+ VDDI VSSI WLP_SAEB_L1 WLP_SAEB_R2 S1AHSF400W40_IO_SIM
XIO_LR AWT2_L2 AWT2_L1 BIST2IO_L2 BIST2IO_L1 BWEBM_LR BWEB_LR CKD_L2 CKD_L1 
+ DM_LR D_LR GBLB_LR_12 GBL_LR_12 GWB_LR_12 GW_LR_12 PD_BUF_L2 PD_BUF_1 Q_LR 
+ VDDHD VDDI VSSI WLP_SAEB_L2 WLP_SAEB_L1 S1AHSF400W40_IO_SIM
XIO_RR AWT2_R3 AWT2_R4 BIST2IO_R3 BIST2IO_R4 NET339 NET334 CKD_R3 CKD_R4 
+ NET333 NET221 NET326 NET324 NET341 NET340 PD_BUF_R3 PD_BUF_R4 NET332 VDDHD 
+ VDDI VSSI WLP_SAEB_R3 WLP_SAEB_R4 S1AHSF400W40_IO_SIM
XTKWL_R VDDI TK_R3 NET415 VSSI WL_DUM_R3 NET408 WL_TK_R3 WL_TK_LD S1AHSF400W40_TKWL_SIM
XTKWL_L VDDI TK TK_R2 VSSI WL_DUM_LT WL_DUM_R2 WL_TK WL_TK_R2 S1AHSF400W40_TKWL_SIM
XTKWL_LD VDDI TK_R2 TK_R3 VSSI WL_DUM_R2 WL_DUM_R3 WL_TK_R2 WL_TK_R3 
+ S1AHSF400W40_TKWL_LD_SIM
XTKBL TRKBL BL_TK_TP VDDHD PD VDDHD VDDI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI WL_TK_ACT[0] 
+ WL_TK_ACT[1] WL_TK_ACT[2] WL_TK_ACT[3] WL_TK_ACT[4] WL_TK_ACT[5] 
+ WL_TK_ACT[6] WL_TK_ACT[7] WL_TK_ACT[8] WL_TK_ACT[9] WL_TK_ACT[10] 
+ WL_TK_ACT[11] WL_TK_ACT[12] WL_TK_ACT[13] WL_TK_ACT[14] WL_TK_ACT[15] 
+ WL_TK_ACT[16] WL_TK_ACT[17] WL_TK_ACT[18] WL_TK_ACT[19] WL_TK_ACT[20] 
+ WL_TK_ACT[21] WL_TK_ACT[22] WL_TK_ACT[23] WL_TK_ACT[24] WL_TK_ACT[25] 
+ WL_TK_ACT[26] WL_TK_ACT[27] WL_TK_ACT[28] WL_TK_ACT[29] WL_TK_ACT[30] 
+ WL_TK_ACT[31] WL_TK_ACT[32] WL_TK_ACT[33] WL_TK_ACT[34] WL_TK_ACT[35] 
+ WL_TK_ACT[36] WL_TK_ACT[37] WL_TK_ACT[38] WL_TK_ACT[39] WL_TK_ACT[40] 
+ WL_TK_ACT[41] WL_TK_ACT[42] WL_TK_ACT[43] WL_TK_ACT[44] WL_TK_ACT[45] 
+ WL_TK_ACT[46] WL_TK_ACT[47] WL_TK_ACT[48] WL_TK_ACT[49] WL_TK_ACT[50] 
+ WL_TK_ACT[51] WL_TK_ACT[52] WL_TK_ACT[53] WL_TK_ACT[54] WL_TK_ACT[55] 
+ WL_TK_ACT[56] WL_TK_ACT[57] WL_TK_ACT[58] WL_TK_ACT[59] WL_TK_ACT[60] 
+ WL_TK_ACT[61] WL_TK_ACT[62] WL_TK_ACT[63] WL_TK_ACT[64] WL_TK_ACT[65] 
+ WL_TK_ACT[66] WL_TK_ACT[67] WL_TK_ACT[68] WL_TK_ACT[69] WL_TK_ACT[70] 
+ WL_TK_ACT[71] WL_TK_ACT[72] WL_TK_ACT[73] WL_TK_ACT[74] WL_TK_ACT[75] 
+ WL_TK_ACT[76] WL_TK_ACT[77] WL_TK_ACT[78] WL_TK_ACT[79] WL_TK_ACT[80] 
+ WL_TK_ACT[81] WL_TK_ACT[82] WL_TK_ACT[83] WL_TK_ACT[84] WL_TK_ACT[85] 
+ WL_TK_ACT[86] WL_TK_ACT[87] WL_TK_ACT[88] WL_TK_ACT[89] WL_TK_ACT[90] 
+ WL_TK_ACT[91] WL_TK_ACT[92] WL_TK_ACT[93] WL_TK_ACT[94] WL_TK_ACT[95] 
+ WL_TK_ACT[96] WL_TK_ACT[97] WL_TK_ACT[98] WL_TK_ACT[99] WL_TK_ACT[100] 
+ WL_TK_ACT[101] WL_TK_ACT[102] WL_TK_ACT[103] WL_TK_ACT[104] WL_TK_ACT[105] 
+ WL_TK_ACT[106] WL_TK_ACT[107] WL_TK_ACT[108] WL_TK_ACT[109] WL_TK_ACT[110] 
+ WL_TK_ACT[111] WL_TK_ACT[112] WL_TK_ACT[113] WL_TK_ACT[114] WL_TK_ACT[115] 
+ WL_TK_ACT[116] WL_TK_ACT[117] WL_TK_ACT[118] WL_TK_ACT[119] WL_TK_ACT[120] 
+ WL_TK_ACT[121] WL_TK_ACT[122] WL_TK_ACT[123] WL_TK_ACT[124] WL_TK_ACT[125] 
+ WL_TK_ACT[126] WL_TK_ACT[127] WL_TK_ACT[128] WL_TK_ACT[129] WL_TK_ACT[130] 
+ WL_TK_ACT[131] WL_TK_ACT[132] WL_TK_ACT[133] WL_TK_ACT[134] WL_TK_ACT[135] 
+ WL_TK_ACT[136] WL_TK_ACT[137] WL_TK_ACT[138] WL_TK_ACT[139] WL_TK_ACT[140] 
+ WL_TK_ACT[141] WL_TK_ACT[142] WL_TK_ACT[143] WL_TK_ACT[144] WL_TK_ACT[145] 
+ WL_TK_ACT[146] WL_TK_ACT[147] WL_TK_ACT[148] WL_TK_ACT[149] WL_TK_ACT[150] 
+ WL_TK_ACT[151] WL_TK_ACT[152] WL_TK_ACT[153] WL_TK_ACT[154] WL_TK_ACT[155] 
+ WL_TK_ACT[156] WL_TK_ACT[157] WL_TK_ACT[158] WL_TK_ACT[159] WL_TK_ACT[160] 
+ WL_TK_ACT[161] WL_TK_ACT[162] WL_TK_ACT[163] WL_TK_ACT[164] WL_TK_ACT[165] 
+ WL_TK_ACT[166] WL_TK_ACT[167] WL_TK_ACT[168] WL_TK_ACT[169] WL_TK_ACT[170] 
+ WL_TK_ACT[171] WL_TK_ACT[172] WL_TK_ACT[173] WL_TK_ACT[174] WL_TK_ACT[175] 
+ WL_TK_ACT[176] WL_TK_ACT[177] WL_TK_ACT[178] WL_TK_ACT[179] WL_TK_ACT[180] 
+ WL_TK_ACT[181] WL_TK_ACT[182] WL_TK_ACT[183] WL_TK_ACT[184] WL_TK_ACT[185] 
+ WL_TK_ACT[186] WL_TK_ACT[187] WL_TK_ACT[188] WL_TK_ACT[189] WL_TK_ACT[190] 
+ WL_TK_ACT[191] WL_TK_ACT[192] WL_TK_ACT[193] WL_TK_ACT[194] WL_TK_ACT[195] 
+ WL_TK_ACT[196] WL_TK_ACT[197] WL_TK_ACT[198] WL_TK_ACT[199] WL_TK_ACT[200] 
+ WL_TK_ACT[201] WL_TK_ACT[202] WL_TK_ACT[203] WL_TK_ACT[204] WL_TK_ACT[205] 
+ WL_TK_ACT[206] WL_TK_ACT[207] WL_TK_ACT[208] WL_TK_ACT[209] WL_TK_ACT[210] 
+ WL_TK_ACT[211] WL_TK_ACT[212] WL_TK_ACT[213] WL_TK_ACT[214] WL_TK_ACT[215] 
+ WL_TK_ACT[216] WL_TK_ACT[217] WL_TK_ACT[218] WL_TK_ACT[219] WL_TK_ACT[220] 
+ WL_TK_ACT[221] WL_TK_ACT[222] WL_TK_ACT[223] WL_TK_ACT[224] WL_TK_ACT[225] 
+ WL_TK_ACT[226] WL_TK_ACT[227] WL_TK_ACT[228] WL_TK_ACT[229] WL_TK_ACT[230] 
+ WL_TK_ACT[231] WL_TK_ACT[232] WL_TK_ACT[233] WL_TK_ACT[234] WL_TK_ACT[235] 
+ WL_TK_ACT[236] WL_TK_ACT[237] WL_TK_ACT[238] WL_TK_ACT[239] WL_TK_ACT[240] 
+ WL_TK_ACT[241] WL_TK_ACT[242] WL_TK_ACT[243] WL_TK_ACT[244] WL_TK_ACT[245] 
+ WL_TK_ACT[246] WL_TK_ACT[247] WL_TK_ACT[248] WL_TK_ACT[249] WL_TK_ACT[250] 
+ WL_TK_ACT[251] WL_TK_ACT[252] WL_TK_ACT[253] WL_TK_ACT[254] WL_TK_ACT[255] 
+ WL_TK_ACT[256] WL_TK_ACT[257] WL_TK_ACT[258] WL_TK_ACT[259] WL_TK_ACT[260] 
+ WL_TK_ACT[261] WL_TK_ACT[262] WL_TK_ACT[263] WL_TK_ACT[264] WL_TK_ACT[265] 
+ WL_TK_ACT[266] WL_TK_ACT[267] WL_TK_ACT[268] WL_TK_ACT[269] WL_TK_ACT[270] 
+ WL_TK_ACT[271] WL_TK_ACT[272] WL_TK_ACT[273] WL_TK_ACT[274] WL_TK_ACT[275] 
+ WL_TK_ACT[276] WL_TK_ACT[277] WL_TK_ACT[278] WL_TK_ACT[279] WL_TK_ACT[280] 
+ WL_TK_ACT[281] WL_TK_ACT[282] WL_TK_ACT[283] WL_TK_ACT[284] WL_TK_ACT[285] 
+ WL_TK_ACT[286] WL_TK_ACT[287] WL_TK_ACT[288] WL_TK_ACT[289] WL_TK_ACT[290] 
+ WL_TK_ACT[291] WL_TK_ACT[292] WL_TK_ACT[293] WL_TK_ACT[294] WL_TK_ACT[295] 
+ WL_TK_ACT[296] WL_TK_ACT[297] WL_TK_ACT[298] WL_TK_ACT[299] WL_TK_ACT[300] 
+ WL_TK_ACT[301] WL_TK_ACT[302] WL_TK_ACT[303] WL_TK_ACT[304] WL_TK_ACT[305] 
+ WL_TK_ACT[306] WL_TK_ACT[307] WL_TK_ACT[308] WL_TK_ACT[309] WL_TK_ACT[310] 
+ WL_TK_ACT[311] WL_TK_ACT[312] WL_TK_ACT[313] WL_TK_ACT[314] WL_TK_ACT[315] 
+ WL_TK_ACT[316] WL_TK_ACT[317] WL_TK_ACT[318] WL_TK_ACT[319] WL_TK_ACT[320] 
+ WL_TK_ACT[321] WL_TK_ACT[322] WL_TK_ACT[323] WL_TK_ACT[324] WL_TK_ACT[325] 
+ WL_TK_ACT[326] WL_TK_ACT[327] WL_TK_ACT[328] WL_TK_ACT[329] WL_TK_ACT[330] 
+ WL_TK_ACT[331] WL_TK_ACT[332] WL_TK_ACT[333] WL_TK_ACT[334] WL_TK_ACT[335] 
+ WL_TK_ACT[336] WL_TK_ACT[337] WL_TK_ACT[338] WL_TK_ACT[339] WL_TK_ACT[340] 
+ WL_TK_ACT[341] WL_TK_ACT[342] WL_TK_ACT[343] WL_TK_ACT[344] WL_TK_ACT[345] 
+ WL_TK_ACT[346] WL_TK_ACT[347] WL_TK_ACT[348] WL_TK_ACT[349] WL_TK_ACT[350] 
+ WL_TK_ACT[351] WL_TK_ACT[352] WL_TK_ACT[353] WL_TK_ACT[354] WL_TK_ACT[355] 
+ WL_TK_ACT[356] WL_TK_ACT[357] WL_TK_ACT[358] WL_TK_ACT[359] WL_TK_ACT[360] 
+ WL_TK_ACT[361] WL_TK_ACT[362] WL_TK_ACT[363] WL_TK_ACT[364] WL_TK_ACT[365] 
+ WL_TK_ACT[366] WL_TK_ACT[367] WL_TK_ACT[368] WL_TK_ACT[369] WL_TK_ACT[370] 
+ WL_TK_ACT[371] WL_TK_ACT[372] WL_TK_ACT[373] WL_TK_ACT[374] WL_TK_ACT[375] 
+ WL_TK_ACT[376] WL_TK_ACT[377] WL_TK_ACT[378] WL_TK_ACT[379] WL_TK_ACT[380] 
+ WL_TK_ACT[381] WL_TK_ACT[382] WL_TK_ACT[383] WL_TK_ACT[384] WL_TK_ACT[385] 
+ WL_TK_ACT[386] WL_TK_ACT[387] WL_TK_ACT[388] WL_TK_ACT[389] WL_TK_ACT[390] 
+ WL_TK_ACT[391] WL_TK_ACT[392] WL_TK_ACT[393] WL_TK_ACT[394] WL_TK_ACT[395] 
+ WL_TK_ACT[396] WL_TK_ACT[397] WL_TK_ACT[398] WL_TK_ACT[399] WL_TK_ACT[400] 
+ WL_TK_ACT[401] WL_TK_ACT[402] WL_TK_ACT[403] WL_TK_ACT[404] WL_TK_ACT[405] 
+ WL_TK_ACT[406] WL_TK_ACT[407] WL_TK_ACT[408] WL_TK_ACT[409] WL_TK_ACT[410] 
+ WL_TK_ACT[411] WL_TK_ACT[412] WL_TK_ACT[413] WL_TK_ACT[414] WL_TK_ACT[415] 
+ WL_TK_ACT[416] WL_TK_ACT[417] WL_TK_ACT[418] WL_TK_ACT[419] WL_TK_ACT[420] 
+ WL_TK_ACT[421] WL_TK_ACT[422] WL_TK_ACT[423] WL_TK_ACT[424] WL_TK_ACT[425] 
+ WL_TK_ACT[426] WL_TK_ACT[427] WL_TK_ACT[428] WL_TK_ACT[429] WL_TK_ACT[430] 
+ WL_TK_ACT[431] WL_TK_ACT[432] WL_TK_ACT[433] WL_TK_ACT[434] WL_TK_ACT[435] 
+ WL_TK_ACT[436] WL_TK_ACT[437] WL_TK_ACT[438] WL_TK_ACT[439] WL_TK_ACT[440] 
+ WL_TK_ACT[441] WL_TK_ACT[442] WL_TK_ACT[443] WL_TK_ACT[444] WL_TK_ACT[445] 
+ WL_TK_ACT[446] WL_TK_ACT[447] WL_TK_ACT[448] WL_TK_ACT[449] WL_TK_ACT[450] 
+ WL_TK_ACT[451] WL_TK_ACT[452] WL_TK_ACT[453] WL_TK_ACT[454] WL_TK_ACT[455] 
+ WL_TK_ACT[456] WL_TK_ACT[457] WL_TK_ACT[458] WL_TK_ACT[459] WL_TK_ACT[460] 
+ WL_TK_ACT[461] WL_TK_ACT[462] WL_TK_ACT[463] WL_TK_ACT[464] WL_TK_ACT[465] 
+ WL_TK_ACT[466] WL_TK_ACT[467] WL_TK_ACT[468] WL_TK_ACT[469] WL_TK_ACT[470] 
+ WL_TK_ACT[471] WL_TK_ACT[472] WL_TK_ACT[473] WL_TK_ACT[474] WL_TK_ACT[475] 
+ WL_TK_ACT[476] WL_TK_ACT[477] WL_TK_ACT[478] WL_TK_ACT[479] WL_TK_ACT[480] 
+ WL_TK_ACT[481] WL_TK_ACT[482] WL_TK_ACT[483] WL_TK_ACT[484] WL_TK_ACT[485] 
+ WL_TK_ACT[486] WL_TK_ACT[487] WL_TK_ACT[488] WL_TK_ACT[489] WL_TK_ACT[490] 
+ WL_TK_ACT[491] WL_TK_ACT[492] WL_TK_ACT[493] WL_TK_ACT[494] WL_TK_ACT[495] 
+ WL_TK_ACT[496] WL_TK_ACT[497] WL_TK_ACT[498] WL_TK_ACT[499] WL_TK_ACT[500] 
+ WL_TK_ACT[501] WL_TK_ACT[502] WL_TK_ACT[503] WL_TK_ACT[504] WL_TK_ACT[505] 
+ WL_TK_ACT[506] WL_TK_ACT[507] WL_TK_ACT[508] WL_TK_ACT[509] WL_TK_ACT[510] 
+ WL_TK_ACT[511] TIEH_BT TIEL S1AHSF400W40_TKBL_SIM
XARRLBLLD_LDL BLB_LL_2 BLB_DUM_LL_2 BLB_LL_3 BLB_DUM_LL_3 BL_LL_2 BL_DUM_LL_2 
+ BL_LL_3 BL_DUM_LL_3 VDDI GBLB_LL_12 GBLB_LL_3 GBL_LL_12 GBL_LL_3 GWB_LL_12 
+ GWB_LL_3 GW_LL_12 GW_LL_3 VDDHD VDDI VSSI S1AHSF400W40_ARR_BLLD_SIM
XARR_BLLD_LDR BLB_LR_2 BLB_DUM_LR_2 BLB_LR_3 BLB_DUM_LR_3 BL_LR_2 BL_DUM_LR_2 
+ BL_LR_3 BL_DUM_LR_3 VDDI GBLB_LR_12 GBLB_LR_3 GBL_LR_12 GBL_LR_3 GWB_LR_12 
+ GWB_LR_3 GW_LR_12 GW_LR_3 VDDHD VDDI VSSI S1AHSF400W40_ARR_BLLD_SIM
XARR_WLLD_LD VDDI VDDHD VDDI VSSI WL_LD3[0] WL_LD3[1] WL_LD2[0] WL_LD2[1] 
+ S1AHSF400W40_ARR_WLLD_SIM
XARR_WLLD_RD VDDI VDDHD VDDI VSSI WL_RD2[0] WL_RD2[1] WL_RD3[0] WL_RD3[1] 
+ S1AHSF400W40_ARR_WLLD_SIM
XARR_MCB_RDR NET0103 NET0100 NET0101 NET0102 VDDI NET098 NET089 NET097 NET099 
+ VDDHD VDDI VSSI WL_RD3[0] WL_RD3[1] WL_RD4[0] WL_RD4[1] S1AHSF400W40_ARR_MCB_SIM
XARR_MCB_RDL NET0113 NET0114 NET0115 NET0112 VDDI NET0116 NET0118 NET0119 
+ NET0117 VDDHD VDDI VSSI WL_RD1[0] WL_RD1[1] WL_RD2[0] WL_RD2[1] S1AHSF400W40_ARR_MCB_SIM
XARR_MCB_LDR BL_LR_2 BL_DUM_LR_2 BLB_LR_2 BLB_DUM_LR_2 VDDI GBL_LR_12 
+ GBLB_LR_12 GW_LR_12 GWB_LR_12 VDDHD VDDI VSSI WL_LD2[0] WL_LD2[1] WL_LD1[0] 
+ WL_LD1[1] S1AHSF400W40_ARR_MCB_SIM
XARR_MCB_LDL BL_LL_2 BL_DUM_LL_2 BLB_LL_2 BLB_DUM_LL_2 VDDI GBL_LL_12 
+ GBLB_LL_12 GW_LL_12 GWB_LL_12 VDDHD VDDI VSSI WL_LD4[0] WL_LD4[1] WL_LD3[0] 
+ WL_LD3[1] S1AHSF400W40_ARR_MCB_SIM
XARR_LIO_RDL NET562 NET0514 NET0513[0] NET0513[1] NET0513[2] NET0513[3] 
+ NET0513[4] NET0513[5] NET0513[6] NET0513[7] NET0513[8] NET0513[9] 
+ NET0513[10] NET0513[11] NET0513[12] NET0513[13] NET580 NET0512 NET0511[0] 
+ NET0511[1] NET0511[2] NET0511[3] NET0511[4] NET0511[5] NET0511[6] NET0511[7] 
+ NET0511[8] NET0511[9] NET0511[10] NET0511[11] NET0511[12] NET0511[13] 
+ BLEQ_DN_RD1 BLEQ_DN_RD2 BLEQ_UP_RD1 BLEQ_UP_RD2 NET150 NET0510 NET0509[0] 
+ NET0509[1] NET0509[2] NET0509[3] NET0509[4] NET0509[5] NET0509[6] NET0509[7] 
+ NET0509[8] NET0509[9] NET0509[10] NET0509[11] NET0509[12] NET0509[13] NET193 
+ NET0508 NET0507[0] NET0507[1] NET0507[2] NET0507[3] NET0507[4] NET0507[5] 
+ NET0507[6] NET0507[7] NET0507[8] NET0507[9] NET0507[10] NET0507[11] 
+ NET0507[12] NET0507[13] VDDI NET147 NET141 NET584 NET583 NET582 NET581 
+ NET189 NET211 RE_RD1 RE_RD2 SAEB_RD1 SAEB_RD2 VDDHD VDDI VSSI WE_RD1 WE_RD2 
+ YL_RD1[0] YL_RD1[1] YL_RD2[0] YL_RD2[1] Y_DN_RD1[0] Y_DN_RD1[1] Y_DN_RD1[2] 
+ Y_DN_RD1[3] Y_DN_RD1[4] Y_DN_RD1[5] Y_DN_RD1[6] Y_DN_RD1[7] Y_DN_RD2[0] 
+ Y_DN_RD2[1] Y_DN_RD2[2] Y_DN_RD2[3] Y_DN_RD2[4] Y_DN_RD2[5] Y_DN_RD2[6] 
+ Y_DN_RD2[7] Y_UP_RD1[0] Y_UP_RD1[1] Y_UP_RD1[2] Y_UP_RD1[3] Y_UP_RD1[4] 
+ Y_UP_RD1[5] Y_UP_RD1[6] Y_UP_RD1[7] Y_UP_RD2[0] Y_UP_RD2[1] Y_UP_RD2[2] 
+ Y_UP_RD2[3] Y_UP_RD2[4] Y_UP_RD2[5] Y_UP_RD2[6] Y_UP_RD2[7] S1AHSF400W40_ARR_LIO_SIM
XARR_LIO_RDR NET598 NET0554 NET0553[0] NET0553[1] NET0553[2] NET0553[3] 
+ NET0553[4] NET0553[5] NET0553[6] NET0553[7] NET0553[8] NET0553[9] 
+ NET0553[10] NET0553[11] NET0553[12] NET0553[13] NET616 NET0552 NET0551[0] 
+ NET0551[1] NET0551[2] NET0551[3] NET0551[4] NET0551[5] NET0551[6] NET0551[7] 
+ NET0551[8] NET0551[9] NET0551[10] NET0551[11] NET0551[12] NET0551[13] 
+ BLEQ_DN_RD3 BLEQ_DN_RD4 BLEQ_UP_RD3 BLEQ_UP_RD4 NET615 NET0550 NET0549[0] 
+ NET0549[1] NET0549[2] NET0549[3] NET0549[4] NET0549[5] NET0549[6] NET0549[7] 
+ NET0549[8] NET0549[9] NET0549[10] NET0549[11] NET0549[12] NET0549[13] NET198 
+ NET0548 NET0547[0] NET0547[1] NET0547[2] NET0547[3] NET0547[4] NET0547[5] 
+ NET0547[6] NET0547[7] NET0547[8] NET0547[9] NET0547[10] NET0547[11] 
+ NET0547[12] NET0547[13] VDDI NET622 NET621 NET620 NET196 NET618 NET617 
+ NET614 NET613 RE_RD3 RE_RD4 SAEB_RD3 SAEB_RD4 VDDHD VDDI VSSI WE_RD3 WE_RD4 
+ YL_RD3[0] YL_RD3[1] YL_RD4[0] YL_RD4[1] Y_DN_RD3[0] Y_DN_RD3[1] Y_DN_RD3[2] 
+ Y_DN_RD3[3] Y_DN_RD3[4] Y_DN_RD3[5] Y_DN_RD3[6] Y_DN_RD3[7] Y_DN_RD4[0] 
+ Y_DN_RD4[1] Y_DN_RD4[2] Y_DN_RD4[3] Y_DN_RD4[4] Y_DN_RD4[5] Y_DN_RD4[6] 
+ Y_DN_RD4[7] Y_UP_RD3[0] Y_UP_RD3[1] Y_UP_RD3[2] Y_UP_RD3[3] Y_UP_RD3[4] 
+ Y_UP_RD3[5] Y_UP_RD3[6] Y_UP_RD3[7] Y_UP_RD4[0] Y_UP_RD4[1] Y_UP_RD4[2] 
+ Y_UP_RD4[3] Y_UP_RD4[4] Y_UP_RD4[5] Y_UP_RD4[6] Y_UP_RD4[7] S1AHSF400W40_ARR_LIO_SIM
XARR_LIO_LDL BLB_LL_3 BLB_DUM_LL_3 NET0593[0] NET0593[1] NET0593[2] NET0593[3] 
+ NET0593[4] NET0593[5] NET0593[6] NET0593[7] NET0593[8] NET0593[9] 
+ NET0593[10] NET0593[11] NET0593[12] NET0593[13] BLB_LL_4 BLB_DUM_LL_4 
+ NET0591[0] NET0591[1] NET0591[2] NET0591[3] NET0591[4] NET0591[5] NET0591[6] 
+ NET0591[7] NET0591[8] NET0591[9] NET0591[10] NET0591[11] NET0591[12] 
+ NET0591[13] BLEQ_DN_LD4 BLEQ_DN_LD3 BLEQ_UP_LD4 BLEQ_UP_LD3 BL_LL_3 
+ BL_DUM_LL_3 NET0589[0] NET0589[1] NET0589[2] NET0589[3] NET0589[4] 
+ NET0589[5] NET0589[6] NET0589[7] NET0589[8] NET0589[9] NET0589[10] 
+ NET0589[11] NET0589[12] NET0589[13] BL_LL_4 BL_DUM_LL_4 NET0587[0] 
+ NET0587[1] NET0587[2] NET0587[3] NET0587[4] NET0587[5] NET0587[6] NET0587[7] 
+ NET0587[8] NET0587[9] NET0587[10] NET0587[11] NET0587[12] NET0587[13] VDDI 
+ GBLB_LL_3 GBLB_LL_4 GBL_LL_3 GBL_LL_4 GWB_LL_3 GWB_LL_4 GW_LL_3 GW_LL_4 
+ RE_LD4 RE_LD3 SAEB_LD4 SAEB_LD3 VDDHD VDDI VSSI WE_LD4 WE_LD3 YL_LD4[0] 
+ YL_LD4[1] YL_LD3[0] YL_LD3[1] Y_DN_LD4[0] Y_DN_LD4[1] Y_DN_LD4[2] 
+ Y_DN_LD4[3] Y_DN_LD4[4] Y_DN_LD4[5] Y_DN_LD4[6] Y_DN_LD4[7] Y_DN_LD3[0] 
+ Y_DN_LD3[1] Y_DN_LD3[2] Y_DN_LD3[3] Y_DN_LD3[4] Y_DN_LD3[5] Y_DN_LD3[6] 
+ Y_DN_LD3[7] Y_UP_LD4[0] Y_UP_LD4[1] Y_UP_LD4[2] Y_UP_LD4[3] Y_UP_LD4[4] 
+ Y_UP_LD4[5] Y_UP_LD4[6] Y_UP_LD4[7] Y_UP_LD3[0] Y_UP_LD3[1] Y_UP_LD3[2] 
+ Y_UP_LD3[3] Y_UP_LD3[4] Y_UP_LD3[5] Y_UP_LD3[6] Y_UP_LD3[7] S1AHSF400W40_ARR_LIO_SIM
XARR_LIO_LDR BLB_LR_3 BLB_DUM_LR_3 NET0633[0] NET0633[1] NET0633[2] NET0633[3] 
+ NET0633[4] NET0633[5] NET0633[6] NET0633[7] NET0633[8] NET0633[9] 
+ NET0633[10] NET0633[11] NET0633[12] NET0633[13] BLB_LR_4 BLB_DUM_LR_4 
+ NET0631[0] NET0631[1] NET0631[2] NET0631[3] NET0631[4] NET0631[5] NET0631[6] 
+ NET0631[7] NET0631[8] NET0631[9] NET0631[10] NET0631[11] NET0631[12] 
+ NET0631[13] BLEQ_DN_LD2 BLEQ_DN_LD1 BLEQ_UP_LD2 BLEQ_UP_LD1 BL_LR_3 
+ BL_DUM_LR_3 NET088[0] NET088[1] NET088[2] NET088[3] NET088[4] NET088[5] 
+ NET088[6] NET088[7] NET088[8] NET088[9] NET088[10] NET088[11] NET088[12] 
+ NET088[13] BL_LR_4 BL_DUM_LR_4 NET0627[0] NET0627[1] NET0627[2] NET0627[3] 
+ NET0627[4] NET0627[5] NET0627[6] NET0627[7] NET0627[8] NET0627[9] 
+ NET0627[10] NET0627[11] NET0627[12] NET0627[13] VDDI GBLB_LR_3 GBLB_LR_4 
+ GBL_LR_3 GBL_LR_4 GWB_LR_3 GWB_LR_4 GW_LR_3 GW_LR_4 RE_LD2 RE_LD1 SAEB_LD2 
+ SAEB_LD1 VDDHD VDDI VSSI WE_LD2 WE_LD1 YL_LD2[0] YL_LD2[1] YL_LD1[0] 
+ YL_LD1[1] Y_DN_LD2[0] Y_DN_LD2[1] Y_DN_LD2[2] Y_DN_LD2[3] Y_DN_LD2[4] 
+ Y_DN_LD2[5] Y_DN_LD2[6] Y_DN_LD2[7] Y_DN_LD1[0] Y_DN_LD1[1] Y_DN_LD1[2] 
+ Y_DN_LD1[3] Y_DN_LD1[4] Y_DN_LD1[5] Y_DN_LD1[6] Y_DN_LD1[7] Y_UP_LD2[0] 
+ Y_UP_LD2[1] Y_UP_LD2[2] Y_UP_LD2[3] Y_UP_LD2[4] Y_UP_LD2[5] Y_UP_LD2[6] 
+ Y_UP_LD2[7] Y_UP_LD1[0] Y_UP_LD1[1] Y_UP_LD1[2] Y_UP_LD1[3] Y_UP_LD1[4] 
+ Y_UP_LD1[5] Y_UP_LD1[6] Y_UP_LD1[7] S1AHSF400W40_ARR_LIO_SIM
XARR_LIO_LD_RD BLEQ_DN_RD2 BLEQ_DN_RD3 BLEQ_UP_RD2 BLEQ_UP_RD3 VDDI RE_RD2 
+ RE_RD3 SAEB_RD2 SAEB_RD3 VDDHD VDDI VSSI WE_RD2 WE_RD3 YL_RD2[0] YL_RD2[1] 
+ YL_RD3[0] YL_RD3[1] Y_DN_RD2[0] Y_DN_RD2[1] Y_DN_RD2[2] Y_DN_RD2[3] 
+ Y_DN_RD2[4] Y_DN_RD2[5] Y_DN_RD2[6] Y_DN_RD2[7] Y_DN_RD3[0] Y_DN_RD3[1] 
+ Y_DN_RD3[2] Y_DN_RD3[3] Y_DN_RD3[4] Y_DN_RD3[5] Y_DN_RD3[6] Y_DN_RD3[7] 
+ Y_UP_RD2[0] Y_UP_RD2[1] Y_UP_RD2[2] Y_UP_RD2[3] Y_UP_RD2[4] Y_UP_RD2[5] 
+ Y_UP_RD2[6] Y_UP_RD2[7] Y_UP_RD3[0] Y_UP_RD3[1] Y_UP_RD3[2] Y_UP_RD3[3] 
+ Y_UP_RD3[4] Y_UP_RD3[5] Y_UP_RD3[6] Y_UP_RD3[7] S1AHSF400W40_ARR_LIO_LD_SIM
XARR_LIO_LD_LD BLEQ_DN_LD3 BLEQ_DN_LD2 BLEQ_UP_LD3 BLEQ_UP_LD2 VDDI RE_LD3 
+ RE_LD2 SAEB_LD3 SAEB_LD2 VDDHD VDDI VSSI WE_LD3 WE_LD2 YL_LD3[0] YL_LD3[1] 
+ YL_LD2[0] YL_LD2[1] Y_DN_LD3[0] Y_DN_LD3[1] Y_DN_LD3[2] Y_DN_LD3[3] 
+ Y_DN_LD3[4] Y_DN_LD3[5] Y_DN_LD3[6] Y_DN_LD3[7] Y_DN_LD2[0] Y_DN_LD2[1] 
+ Y_DN_LD2[2] Y_DN_LD2[3] Y_DN_LD2[4] Y_DN_LD2[5] Y_DN_LD2[6] Y_DN_LD2[7] 
+ Y_UP_LD3[0] Y_UP_LD3[1] Y_UP_LD3[2] Y_UP_LD3[3] Y_UP_LD3[4] Y_UP_LD3[5] 
+ Y_UP_LD3[6] Y_UP_LD3[7] Y_UP_LD2[0] Y_UP_LD2[1] Y_UP_LD2[2] Y_UP_LD2[3] 
+ Y_UP_LD2[4] Y_UP_LD2[5] Y_UP_LD2[6] Y_UP_LD2[7] S1AHSF400W40_ARR_LIO_LD_SIM
XBK_TOP_EDGE VDDHD VDDI VSSI WLP_SAE_4 WLP_SAE_TK_4 S1AHSF400W40_BK_TOP_EDGE_SIM
XTRKPRE PD TRKBL WL_TK VDDHD VDDI VSSI TIEH_BT TIEL S1AHSF400W40_TRKPRE_SIM
XBK_WLDV_LD_D VDDHD VDDI DEC_X0_2[0] DEC_X0_2[1] DEC_X0_2[2] DEC_X0_2[3] 
+ DEC_X0_2[4] DEC_X0_2[5] DEC_X0_2[6] DEC_X0_2[7] DEC_X0_3[0] DEC_X0_3[1] 
+ DEC_X0_3[2] DEC_X0_3[3] DEC_X0_3[4] DEC_X0_3[5] DEC_X0_3[6] DEC_X0_3[7] 
+ DEC_X1_2[0] DEC_X1_2[1] DEC_X1_2[2] DEC_X1_2[3] DEC_X1_2[4] DEC_X1_2[5] 
+ DEC_X1_2[6] DEC_X1_2[7] DEC_X1_3[0] DEC_X1_3[1] DEC_X1_3[2] DEC_X1_3[3] 
+ DEC_X1_3[4] DEC_X1_3[5] DEC_X1_3[6] DEC_X1_3[7] DEC_X2_2[0] DEC_X2_2[1] 
+ DEC_X2_2[2] DEC_X2_2[3] DEC_X2_3[0] DEC_X2_3[1] DEC_X2_3[2] DEC_X2_3[3] 
+ DEC_X3_2[0] DEC_X3_2[1] DEC_X3_2[2] DEC_X3_2[3] DEC_X3_2[4] DEC_X3_2[5] 
+ DEC_X3_2[6] DEC_X3_2[7] DEC_X3_3[0] DEC_X3_3[1] DEC_X3_3[2] DEC_X3_3[3] 
+ DEC_X3_3[4] DEC_X3_3[5] DEC_X3_3[6] DEC_X3_3[7] DEC_Y_2[0] DEC_Y_2[1] 
+ DEC_Y_2[2] DEC_Y_2[3] DEC_Y_2[4] DEC_Y_2[5] DEC_Y_2[6] DEC_Y_2[7] DEC_Y_3[0] 
+ DEC_Y_3[1] DEC_Y_3[2] DEC_Y_3[3] DEC_Y_3[4] DEC_Y_3[5] DEC_Y_3[6] DEC_Y_3[7] 
+ PD_BUF_2 PD_BUF_3 PD_CVDDBUF_2 PD_CVDDBUF_3 RW_RE_2 RW_RE_3 VDDHD VDDI VSSI 
+ WLP_SAE_2 WLP_SAE_TK_2 WLP_SAE_TK_3 WLP_SAE_3 YL_2[0] YL_3[0] 
+ S1AHSF400W40_BK_WLDV_LD_SIM
XBK_LCNT_D BLEQ_DN_LD1 BLEQ_DN_RD1 BLEQ_UP_LD1 BLEQ_UP_RD1 VDDHD VDDI 
+ DEC_X0_3[0] DEC_X0_3[1] DEC_X0_3[2] DEC_X0_3[3] DEC_X0_3[4] DEC_X0_3[5] 
+ DEC_X0_3[6] DEC_X0_3[7] NET0827[0] NET0827[1] NET0827[2] NET0827[3] 
+ NET0827[4] NET0827[5] NET0827[6] NET0827[7] DEC_X1_3[0] DEC_X1_3[1] 
+ DEC_X1_3[2] DEC_X1_3[3] DEC_X1_3[4] DEC_X1_3[5] DEC_X1_3[6] DEC_X1_3[7] 
+ NET0826[0] NET0826[1] NET0826[2] NET0826[3] NET0826[4] NET0826[5] NET0826[6] 
+ NET0826[7] DEC_X2_3[0] DEC_X2_3[1] DEC_X2_3[2] DEC_X2_3[3] NET0824[0] 
+ NET0824[1] NET0824[2] NET0824[3] DEC_X3_3[0] DEC_X3_3[1] DEC_X3_3[2] 
+ DEC_X3_3[3] DEC_X3_3[4] DEC_X3_3[5] DEC_X3_3[6] DEC_X3_3[7] NET0832[0] 
+ NET0832[1] NET0832[2] NET0832[3] NET0832[4] NET0832[5] NET0832[6] NET0832[7] 
+ DEC_Y_3[0] DEC_Y_3[1] DEC_Y_3[2] DEC_Y_3[3] DEC_Y_3[4] DEC_Y_3[5] DEC_Y_3[6] 
+ DEC_Y_3[7] Y_DN_LD1[0] Y_DN_LD1[1] Y_DN_LD1[2] Y_DN_LD1[3] Y_DN_LD1[4] 
+ Y_DN_LD1[5] Y_DN_LD1[6] Y_DN_LD1[7] Y_DN_RD1[0] Y_DN_RD1[1] Y_DN_RD1[2] 
+ Y_DN_RD1[3] Y_DN_RD1[4] Y_DN_RD1[5] Y_DN_RD1[6] Y_DN_RD1[7] NET093[0] 
+ NET093[1] NET093[2] NET093[3] NET093[4] NET093[5] NET093[6] NET093[7] 
+ Y_UP_LD1[0] Y_UP_LD1[1] Y_UP_LD1[2] Y_UP_LD1[3] Y_UP_LD1[4] Y_UP_LD1[5] 
+ Y_UP_LD1[6] Y_UP_LD1[7] Y_UP_RD1[0] Y_UP_RD1[1] Y_UP_RD1[2] Y_UP_RD1[3] 
+ Y_UP_RD1[4] Y_UP_RD1[5] Y_UP_RD1[6] Y_UP_RD1[7] PD_BUF_3 NET095 PD_CVDDBUF_3 
+ NET0840 RE_LD1 RE_RD1 RW_RE_3 NET0842 SAEB_LD1 SAEB_RD1 VDDHD VDDI VSSI 
+ WE_LD1 WE_RD1 WLPYB_3 NET047 WLPY_3 NET0811 WLP_SAE_3 WLP_SAE_TK_3 
+ WLP_SAE_TK_4 WLP_SAE_4 YL_3[0] YL_LD1[0] YL_LD1[1] YL_RD1[0] YL_RD1[1] 
+ NET0825 S1AHSF400W40_BK_LCNT_D_SIM
XWLPY_LD_D VDDHD VDDI VDDHD VDDI VSSI WLPYB_2 WLPYB_3 WLPY_2 WLPY_3 
+ S1AHSF400W40_WLPY_LD_SIM
XBK_WLDV_D VDDHD VDDI DEC_X0_1[0] DEC_X0_1[1] DEC_X0_1[2] DEC_X0_1[3] 
+ DEC_X0_1[4] DEC_X0_1[5] DEC_X0_1[6] DEC_X0_1[7] DEC_X0_2[0] DEC_X0_2[1] 
+ DEC_X0_2[2] DEC_X0_2[3] DEC_X0_2[4] DEC_X0_2[5] DEC_X0_2[6] DEC_X0_2[7] 
+ DEC_X1_1[0] DEC_X1_1[1] DEC_X1_1[2] DEC_X1_1[3] DEC_X1_1[4] DEC_X1_1[5] 
+ DEC_X1_1[6] DEC_X1_1[7] DEC_X1_2[0] DEC_X1_2[1] DEC_X1_2[2] DEC_X1_2[3] 
+ DEC_X1_2[4] DEC_X1_2[5] DEC_X1_2[6] DEC_X1_2[7] DEC_X2_1[0] DEC_X2_1[1] 
+ DEC_X2_1[2] DEC_X2_1[3] DEC_X2_2[0] DEC_X2_2[1] DEC_X2_2[2] DEC_X2_2[3] 
+ DEC_X3_1[0] DEC_X3_1[1] DEC_X3_1[2] DEC_X3_1[3] DEC_X3_1[4] DEC_X3_1[5] 
+ DEC_X3_1[6] DEC_X3_1[7] DEC_X3_2[0] DEC_X3_2[1] DEC_X3_2[2] DEC_X3_2[3] 
+ DEC_X3_2[4] DEC_X3_2[5] DEC_X3_2[6] DEC_X3_2[7] DEC_Y_1[0] DEC_Y_1[1] 
+ DEC_Y_1[2] DEC_Y_1[3] DEC_Y_1[4] DEC_Y_1[5] DEC_Y_1[6] DEC_Y_1[7] DEC_Y_2[0] 
+ DEC_Y_2[1] DEC_Y_2[2] DEC_Y_2[3] DEC_Y_2[4] DEC_Y_2[5] DEC_Y_2[6] DEC_Y_2[7] 
+ PD_BUF_1 PD_BUF_2 PD_CVDDBUF_1 PD_CVDDBUF_2 RW_RE_1 RW_RE_2 VDDHD VDDI VSSI 
+ NET821 WLPYB_2 NET826 WLPY_2 WLP_SAE_1 WLP_SAE_TK_1 WLP_SAE_TK_2 WLP_SAE_2 
+ WL_LD1[0] WL_LD1[1] WL_RD1[0] WL_RD1[1] YL_1[0] YL_2[0] S1AHSF400W40_BK_WLDV_D_SIM
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_WLDV_U
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_WLDV_U DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] 
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] 
+ DEC_Y[7] PD_BUF RW_RE VDDHD VDDI VSSI WL[0] WL[1] WLPY WLPYB WLP_SAE 
+ WLP_SAE_TK YL[0]
*.PININFO WL[0]:O WL[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B PD_BUF:B RW_RE:B VDDHD:B VDDI:B VSSI:B WLPY:B WLPYB:B 
*.PININFO WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XWLDV_0 DEC_X0[6] DEC_X0[7] NET046[0] NET046[1] NET046[2] NET046[3] NET046[4] 
+ NET046[5] DEC_X1[7] NET044[0] NET044[1] NET044[2] NET044[3] NET044[4] 
+ NET044[5] NET044[6] NET040[0] NET040[1] NET040[2] NET040[3] NET041[0] 
+ NET041[1] NET041[2] NET041[3] NET041[4] NET041[5] NET041[6] NET041[7] 
+ NET043[0] NET043[1] NET043[2] NET043[3] NET043[4] NET043[5] NET043[6] 
+ NET043[7] PD_BUF NET29 NET039 VDDHD VDDI VSSI WL[0] WL[1] WLPY WLPYB NET038 
+ NET014 NET042 S1AHSF400W40_XDRV_LA512
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_WLDV_U_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_WLDV_U_SIM CVDDHD CVDDI DEC_X0_BT[0] DEC_X0_BT[1] DEC_X0_BT[2] 
+ DEC_X0_BT[3] DEC_X0_BT[4] DEC_X0_BT[5] DEC_X0_BT[6] DEC_X0_BT[7] 
+ DEC_X0_TP[0] DEC_X0_TP[1] DEC_X0_TP[2] DEC_X0_TP[3] DEC_X0_TP[4] 
+ DEC_X0_TP[5] DEC_X0_TP[6] DEC_X0_TP[7] DEC_X1_BT[0] DEC_X1_BT[1] 
+ DEC_X1_BT[2] DEC_X1_BT[3] DEC_X1_BT[4] DEC_X1_BT[5] DEC_X1_BT[6] 
+ DEC_X1_BT[7] DEC_X1_TP[0] DEC_X1_TP[1] DEC_X1_TP[2] DEC_X1_TP[3] 
+ DEC_X1_TP[4] DEC_X1_TP[5] DEC_X1_TP[6] DEC_X1_TP[7] DEC_X2_BT[0] 
+ DEC_X2_BT[1] DEC_X2_BT[2] DEC_X2_BT[3] DEC_X2_TP[0] DEC_X2_TP[1] 
+ DEC_X2_TP[2] DEC_X2_TP[3] DEC_X3_BT[0] DEC_X3_BT[1] DEC_X3_BT[2] 
+ DEC_X3_BT[3] DEC_X3_BT[4] DEC_X3_BT[5] DEC_X3_BT[6] DEC_X3_BT[7] 
+ DEC_X3_TP[0] DEC_X3_TP[1] DEC_X3_TP[2] DEC_X3_TP[3] DEC_X3_TP[4] 
+ DEC_X3_TP[5] DEC_X3_TP[6] DEC_X3_TP[7] DEC_Y_BT[0] DEC_Y_BT[1] DEC_Y_BT[2] 
+ DEC_Y_BT[3] DEC_Y_BT[4] DEC_Y_BT[5] DEC_Y_BT[6] DEC_Y_BT[7] DEC_Y_TP[0] 
+ DEC_Y_TP[1] DEC_Y_TP[2] DEC_Y_TP[3] DEC_Y_TP[4] DEC_Y_TP[5] DEC_Y_TP[6] 
+ DEC_Y_TP[7] PD_BUF_BT PD_BUF_TP PD_CVDDBUF_BT PD_CVDDBUF_TP RW_RE_BT 
+ RW_RE_TP VDDHD VDDI VSSI WLPYB_BT WLPYB_TP WLPY_BT WLPY_TP WLP_SAE_BT 
+ WLP_SAE_TK_BT WLP_SAE_TK_TP WLP_SAE_TP WL_LT[0] WL_LT[1] WL_RT[0] WL_RT[1] 
+ YL_BT[0] YL_TP[0]
*.PININFO DEC_X0_BT[0]:I DEC_X0_BT[1]:I DEC_X0_BT[2]:I DEC_X0_BT[3]:I 
*.PININFO DEC_X0_BT[4]:I DEC_X0_BT[5]:I DEC_X0_BT[6]:I DEC_X0_BT[7]:I 
*.PININFO DEC_X1_BT[0]:I DEC_X1_BT[1]:I DEC_X1_BT[2]:I DEC_X1_BT[3]:I 
*.PININFO DEC_X1_BT[4]:I DEC_X1_BT[5]:I DEC_X1_BT[6]:I DEC_X1_BT[7]:I 
*.PININFO PD_BUF_BT:I PD_CVDDBUF_BT:I RW_RE_TP:I DEC_X0_TP[0]:O DEC_X0_TP[1]:O 
*.PININFO DEC_X0_TP[2]:O DEC_X0_TP[3]:O DEC_X0_TP[4]:O DEC_X0_TP[5]:O 
*.PININFO DEC_X0_TP[6]:O DEC_X0_TP[7]:O DEC_X1_TP[0]:O DEC_X1_TP[1]:O 
*.PININFO DEC_X1_TP[2]:O DEC_X1_TP[3]:O DEC_X1_TP[4]:O DEC_X1_TP[5]:O 
*.PININFO DEC_X1_TP[6]:O DEC_X1_TP[7]:O PD_BUF_TP:O PD_CVDDBUF_TP:O CVDDHD:B 
*.PININFO CVDDI:B DEC_X2_BT[0]:B DEC_X2_BT[1]:B DEC_X2_BT[2]:B DEC_X2_BT[3]:B 
*.PININFO DEC_X2_TP[0]:B DEC_X2_TP[1]:B DEC_X2_TP[2]:B DEC_X2_TP[3]:B 
*.PININFO DEC_X3_BT[0]:B DEC_X3_BT[1]:B DEC_X3_BT[2]:B DEC_X3_BT[3]:B 
*.PININFO DEC_X3_BT[4]:B DEC_X3_BT[5]:B DEC_X3_BT[6]:B DEC_X3_BT[7]:B 
*.PININFO DEC_X3_TP[0]:B DEC_X3_TP[1]:B DEC_X3_TP[2]:B DEC_X3_TP[3]:B 
*.PININFO DEC_X3_TP[4]:B DEC_X3_TP[5]:B DEC_X3_TP[6]:B DEC_X3_TP[7]:B 
*.PININFO DEC_Y_BT[0]:B DEC_Y_BT[1]:B DEC_Y_BT[2]:B DEC_Y_BT[3]:B 
*.PININFO DEC_Y_BT[4]:B DEC_Y_BT[5]:B DEC_Y_BT[6]:B DEC_Y_BT[7]:B 
*.PININFO DEC_Y_TP[0]:B DEC_Y_TP[1]:B DEC_Y_TP[2]:B DEC_Y_TP[3]:B 
*.PININFO DEC_Y_TP[4]:B DEC_Y_TP[5]:B DEC_Y_TP[6]:B DEC_Y_TP[7]:B RW_RE_BT:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLPYB_BT:B WLPYB_TP:B WLPY_BT:B WLPY_TP:B 
*.PININFO WLP_SAE_BT:B WLP_SAE_TK_BT:B WLP_SAE_TK_TP:B WLP_SAE_TP:B WL_LT[0]:B 
*.PININFO WL_LT[1]:B WL_RT[0]:B WL_RT[1]:B YL_BT[0]:B YL_TP[0]:B
XI24 NET038[0] NET038[1] NET038[2] NET038[3] NET038[4] NET038[5] NET038[6] 
+ NET038[7] NET037[0] NET037[1] NET037[2] NET037[3] NET037[4] NET037[5] 
+ NET037[6] NET037[7] NET036[0] NET036[1] NET036[2] NET036[3] NET035[0] 
+ NET035[1] NET035[2] NET035[3] NET035[4] NET035[5] NET035[6] NET035[7] 
+ NET034[0] NET034[1] NET034[2] NET034[3] NET034[4] NET034[5] NET034[6] 
+ NET034[7] NET31 NET033 NET38 NET32 NET37 NET34[0] NET34[1] NET33 NET30 
+ NET032 NET031 NET03 S1AHSF400W40_BK_WLDV_U
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SIM_1B
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SIM_1B AWT BIST BWEBM_LL BWEBM_LR BWEB_LL BWEB_LR CEB CEBM CLK DM_LL 
+ DM_LR D_LL D_LR FAD1[0] FAD1[1] FAD1[2] FAD1[3] FAD1[4] FAD1[5] FAD1[6] 
+ FAD1[7] FAD1[8] FAD1[9] FAD1[10] FAD2[0] FAD2[1] FAD2[2] FAD2[3] FAD2[4] 
+ FAD2[5] FAD2[6] FAD2[7] FAD2[8] FAD2[9] FAD2[10] PD PTSEL Q_LL Q_LR REDEN1 
+ REDEN2 RSTB RTSEL[0] RTSEL[1] SCLK SDIN SDOUT TM VDDI VSSI WEB WEBM 
+ WL_TK_ACT[0] WL_TK_ACT[1] WL_TK_ACT[2] WL_TK_ACT[3] WL_TK_ACT[4] 
+ WL_TK_ACT[5] WL_TK_ACT[6] WL_TK_ACT[7] WL_TK_ACT[8] WL_TK_ACT[9] 
+ WL_TK_ACT[10] WL_TK_ACT[11] WL_TK_ACT[12] WL_TK_ACT[13] WL_TK_ACT[14] 
+ WL_TK_ACT[15] WL_TK_ACT[16] WL_TK_ACT[17] WL_TK_ACT[18] WL_TK_ACT[19] 
+ WL_TK_ACT[20] WL_TK_ACT[21] WL_TK_ACT[22] WL_TK_ACT[23] WL_TK_ACT[24] 
+ WL_TK_ACT[25] WL_TK_ACT[26] WL_TK_ACT[27] WL_TK_ACT[28] WL_TK_ACT[29] 
+ WL_TK_ACT[30] WL_TK_ACT[31] WL_TK_ACT[32] WL_TK_ACT[33] WL_TK_ACT[34] 
+ WL_TK_ACT[35] WL_TK_ACT[36] WL_TK_ACT[37] WL_TK_ACT[38] WL_TK_ACT[39] 
+ WL_TK_ACT[40] WL_TK_ACT[41] WL_TK_ACT[42] WL_TK_ACT[43] WL_TK_ACT[44] 
+ WL_TK_ACT[45] WL_TK_ACT[46] WL_TK_ACT[47] WL_TK_ACT[48] WL_TK_ACT[49] 
+ WL_TK_ACT[50] WL_TK_ACT[51] WL_TK_ACT[52] WL_TK_ACT[53] WL_TK_ACT[54] 
+ WL_TK_ACT[55] WL_TK_ACT[56] WL_TK_ACT[57] WL_TK_ACT[58] WL_TK_ACT[59] 
+ WL_TK_ACT[60] WL_TK_ACT[61] WL_TK_ACT[62] WL_TK_ACT[63] WL_TK_ACT[64] 
+ WL_TK_ACT[65] WL_TK_ACT[66] WL_TK_ACT[67] WL_TK_ACT[68] WL_TK_ACT[69] 
+ WL_TK_ACT[70] WL_TK_ACT[71] WL_TK_ACT[72] WL_TK_ACT[73] WL_TK_ACT[74] 
+ WL_TK_ACT[75] WL_TK_ACT[76] WL_TK_ACT[77] WL_TK_ACT[78] WL_TK_ACT[79] 
+ WL_TK_ACT[80] WL_TK_ACT[81] WL_TK_ACT[82] WL_TK_ACT[83] WL_TK_ACT[84] 
+ WL_TK_ACT[85] WL_TK_ACT[86] WL_TK_ACT[87] WL_TK_ACT[88] WL_TK_ACT[89] 
+ WL_TK_ACT[90] WL_TK_ACT[91] WL_TK_ACT[92] WL_TK_ACT[93] WL_TK_ACT[94] 
+ WL_TK_ACT[95] WL_TK_ACT[96] WL_TK_ACT[97] WL_TK_ACT[98] WL_TK_ACT[99] 
+ WL_TK_ACT[100] WL_TK_ACT[101] WL_TK_ACT[102] WL_TK_ACT[103] WL_TK_ACT[104] 
+ WL_TK_ACT[105] WL_TK_ACT[106] WL_TK_ACT[107] WL_TK_ACT[108] WL_TK_ACT[109] 
+ WL_TK_ACT[110] WL_TK_ACT[111] WL_TK_ACT[112] WL_TK_ACT[113] WL_TK_ACT[114] 
+ WL_TK_ACT[115] WL_TK_ACT[116] WL_TK_ACT[117] WL_TK_ACT[118] WL_TK_ACT[119] 
+ WL_TK_ACT[120] WL_TK_ACT[121] WL_TK_ACT[122] WL_TK_ACT[123] WL_TK_ACT[124] 
+ WL_TK_ACT[125] WL_TK_ACT[126] WL_TK_ACT[127] WL_TK_ACT[128] WL_TK_ACT[129] 
+ WL_TK_ACT[130] WL_TK_ACT[131] WL_TK_ACT[132] WL_TK_ACT[133] WL_TK_ACT[134] 
+ WL_TK_ACT[135] WL_TK_ACT[136] WL_TK_ACT[137] WL_TK_ACT[138] WL_TK_ACT[139] 
+ WL_TK_ACT[140] WL_TK_ACT[141] WL_TK_ACT[142] WL_TK_ACT[143] WL_TK_ACT[144] 
+ WL_TK_ACT[145] WL_TK_ACT[146] WL_TK_ACT[147] WL_TK_ACT[148] WL_TK_ACT[149] 
+ WL_TK_ACT[150] WL_TK_ACT[151] WL_TK_ACT[152] WL_TK_ACT[153] WL_TK_ACT[154] 
+ WL_TK_ACT[155] WL_TK_ACT[156] WL_TK_ACT[157] WL_TK_ACT[158] WL_TK_ACT[159] 
+ WL_TK_ACT[160] WL_TK_ACT[161] WL_TK_ACT[162] WL_TK_ACT[163] WL_TK_ACT[164] 
+ WL_TK_ACT[165] WL_TK_ACT[166] WL_TK_ACT[167] WL_TK_ACT[168] WL_TK_ACT[169] 
+ WL_TK_ACT[170] WL_TK_ACT[171] WL_TK_ACT[172] WL_TK_ACT[173] WL_TK_ACT[174] 
+ WL_TK_ACT[175] WL_TK_ACT[176] WL_TK_ACT[177] WL_TK_ACT[178] WL_TK_ACT[179] 
+ WL_TK_ACT[180] WL_TK_ACT[181] WL_TK_ACT[182] WL_TK_ACT[183] WL_TK_ACT[184] 
+ WL_TK_ACT[185] WL_TK_ACT[186] WL_TK_ACT[187] WL_TK_ACT[188] WL_TK_ACT[189] 
+ WL_TK_ACT[190] WL_TK_ACT[191] WL_TK_ACT[192] WL_TK_ACT[193] WL_TK_ACT[194] 
+ WL_TK_ACT[195] WL_TK_ACT[196] WL_TK_ACT[197] WL_TK_ACT[198] WL_TK_ACT[199] 
+ WL_TK_ACT[200] WL_TK_ACT[201] WL_TK_ACT[202] WL_TK_ACT[203] WL_TK_ACT[204] 
+ WL_TK_ACT[205] WL_TK_ACT[206] WL_TK_ACT[207] WL_TK_ACT[208] WL_TK_ACT[209] 
+ WL_TK_ACT[210] WL_TK_ACT[211] WL_TK_ACT[212] WL_TK_ACT[213] WL_TK_ACT[214] 
+ WL_TK_ACT[215] WL_TK_ACT[216] WL_TK_ACT[217] WL_TK_ACT[218] WL_TK_ACT[219] 
+ WL_TK_ACT[220] WL_TK_ACT[221] WL_TK_ACT[222] WL_TK_ACT[223] WL_TK_ACT[224] 
+ WL_TK_ACT[225] WL_TK_ACT[226] WL_TK_ACT[227] WL_TK_ACT[228] WL_TK_ACT[229] 
+ WL_TK_ACT[230] WL_TK_ACT[231] WL_TK_ACT[232] WL_TK_ACT[233] WL_TK_ACT[234] 
+ WL_TK_ACT[235] WL_TK_ACT[236] WL_TK_ACT[237] WL_TK_ACT[238] WL_TK_ACT[239] 
+ WL_TK_ACT[240] WL_TK_ACT[241] WL_TK_ACT[242] WL_TK_ACT[243] WL_TK_ACT[244] 
+ WL_TK_ACT[245] WL_TK_ACT[246] WL_TK_ACT[247] WL_TK_ACT[248] WL_TK_ACT[249] 
+ WL_TK_ACT[250] WL_TK_ACT[251] WL_TK_ACT[252] WL_TK_ACT[253] WL_TK_ACT[254] 
+ WL_TK_ACT[255] WL_TK_ACT[256] WL_TK_ACT[257] WL_TK_ACT[258] WL_TK_ACT[259] 
+ WL_TK_ACT[260] WL_TK_ACT[261] WL_TK_ACT[262] WL_TK_ACT[263] WL_TK_ACT[264] 
+ WL_TK_ACT[265] WL_TK_ACT[266] WL_TK_ACT[267] WL_TK_ACT[268] WL_TK_ACT[269] 
+ WL_TK_ACT[270] WL_TK_ACT[271] WL_TK_ACT[272] WL_TK_ACT[273] WL_TK_ACT[274] 
+ WL_TK_ACT[275] WL_TK_ACT[276] WL_TK_ACT[277] WL_TK_ACT[278] WL_TK_ACT[279] 
+ WL_TK_ACT[280] WL_TK_ACT[281] WL_TK_ACT[282] WL_TK_ACT[283] WL_TK_ACT[284] 
+ WL_TK_ACT[285] WL_TK_ACT[286] WL_TK_ACT[287] WL_TK_ACT[288] WL_TK_ACT[289] 
+ WL_TK_ACT[290] WL_TK_ACT[291] WL_TK_ACT[292] WL_TK_ACT[293] WL_TK_ACT[294] 
+ WL_TK_ACT[295] WL_TK_ACT[296] WL_TK_ACT[297] WL_TK_ACT[298] WL_TK_ACT[299] 
+ WL_TK_ACT[300] WL_TK_ACT[301] WL_TK_ACT[302] WL_TK_ACT[303] WL_TK_ACT[304] 
+ WL_TK_ACT[305] WL_TK_ACT[306] WL_TK_ACT[307] WL_TK_ACT[308] WL_TK_ACT[309] 
+ WL_TK_ACT[310] WL_TK_ACT[311] WL_TK_ACT[312] WL_TK_ACT[313] WL_TK_ACT[314] 
+ WL_TK_ACT[315] WL_TK_ACT[316] WL_TK_ACT[317] WL_TK_ACT[318] WL_TK_ACT[319] 
+ WL_TK_ACT[320] WL_TK_ACT[321] WL_TK_ACT[322] WL_TK_ACT[323] WL_TK_ACT[324] 
+ WL_TK_ACT[325] WL_TK_ACT[326] WL_TK_ACT[327] WL_TK_ACT[328] WL_TK_ACT[329] 
+ WL_TK_ACT[330] WL_TK_ACT[331] WL_TK_ACT[332] WL_TK_ACT[333] WL_TK_ACT[334] 
+ WL_TK_ACT[335] WL_TK_ACT[336] WL_TK_ACT[337] WL_TK_ACT[338] WL_TK_ACT[339] 
+ WL_TK_ACT[340] WL_TK_ACT[341] WL_TK_ACT[342] WL_TK_ACT[343] WL_TK_ACT[344] 
+ WL_TK_ACT[345] WL_TK_ACT[346] WL_TK_ACT[347] WL_TK_ACT[348] WL_TK_ACT[349] 
+ WL_TK_ACT[350] WL_TK_ACT[351] WL_TK_ACT[352] WL_TK_ACT[353] WL_TK_ACT[354] 
+ WL_TK_ACT[355] WL_TK_ACT[356] WL_TK_ACT[357] WL_TK_ACT[358] WL_TK_ACT[359] 
+ WL_TK_ACT[360] WL_TK_ACT[361] WL_TK_ACT[362] WL_TK_ACT[363] WL_TK_ACT[364] 
+ WL_TK_ACT[365] WL_TK_ACT[366] WL_TK_ACT[367] WL_TK_ACT[368] WL_TK_ACT[369] 
+ WL_TK_ACT[370] WL_TK_ACT[371] WL_TK_ACT[372] WL_TK_ACT[373] WL_TK_ACT[374] 
+ WL_TK_ACT[375] WL_TK_ACT[376] WL_TK_ACT[377] WL_TK_ACT[378] WL_TK_ACT[379] 
+ WL_TK_ACT[380] WL_TK_ACT[381] WL_TK_ACT[382] WL_TK_ACT[383] WL_TK_ACT[384] 
+ WL_TK_ACT[385] WL_TK_ACT[386] WL_TK_ACT[387] WL_TK_ACT[388] WL_TK_ACT[389] 
+ WL_TK_ACT[390] WL_TK_ACT[391] WL_TK_ACT[392] WL_TK_ACT[393] WL_TK_ACT[394] 
+ WL_TK_ACT[395] WL_TK_ACT[396] WL_TK_ACT[397] WL_TK_ACT[398] WL_TK_ACT[399] 
+ WL_TK_ACT[400] WL_TK_ACT[401] WL_TK_ACT[402] WL_TK_ACT[403] WL_TK_ACT[404] 
+ WL_TK_ACT[405] WL_TK_ACT[406] WL_TK_ACT[407] WL_TK_ACT[408] WL_TK_ACT[409] 
+ WL_TK_ACT[410] WL_TK_ACT[411] WL_TK_ACT[412] WL_TK_ACT[413] WL_TK_ACT[414] 
+ WL_TK_ACT[415] WL_TK_ACT[416] WL_TK_ACT[417] WL_TK_ACT[418] WL_TK_ACT[419] 
+ WL_TK_ACT[420] WL_TK_ACT[421] WL_TK_ACT[422] WL_TK_ACT[423] WL_TK_ACT[424] 
+ WL_TK_ACT[425] WL_TK_ACT[426] WL_TK_ACT[427] WL_TK_ACT[428] WL_TK_ACT[429] 
+ WL_TK_ACT[430] WL_TK_ACT[431] WL_TK_ACT[432] WL_TK_ACT[433] WL_TK_ACT[434] 
+ WL_TK_ACT[435] WL_TK_ACT[436] WL_TK_ACT[437] WL_TK_ACT[438] WL_TK_ACT[439] 
+ WL_TK_ACT[440] WL_TK_ACT[441] WL_TK_ACT[442] WL_TK_ACT[443] WL_TK_ACT[444] 
+ WL_TK_ACT[445] WL_TK_ACT[446] WL_TK_ACT[447] WL_TK_ACT[448] WL_TK_ACT[449] 
+ WL_TK_ACT[450] WL_TK_ACT[451] WL_TK_ACT[452] WL_TK_ACT[453] WL_TK_ACT[454] 
+ WL_TK_ACT[455] WL_TK_ACT[456] WL_TK_ACT[457] WL_TK_ACT[458] WL_TK_ACT[459] 
+ WL_TK_ACT[460] WL_TK_ACT[461] WL_TK_ACT[462] WL_TK_ACT[463] WL_TK_ACT[464] 
+ WL_TK_ACT[465] WL_TK_ACT[466] WL_TK_ACT[467] WL_TK_ACT[468] WL_TK_ACT[469] 
+ WL_TK_ACT[470] WL_TK_ACT[471] WL_TK_ACT[472] WL_TK_ACT[473] WL_TK_ACT[474] 
+ WL_TK_ACT[475] WL_TK_ACT[476] WL_TK_ACT[477] WL_TK_ACT[478] WL_TK_ACT[479] 
+ WL_TK_ACT[480] WL_TK_ACT[481] WL_TK_ACT[482] WL_TK_ACT[483] WL_TK_ACT[484] 
+ WL_TK_ACT[485] WL_TK_ACT[486] WL_TK_ACT[487] WL_TK_ACT[488] WL_TK_ACT[489] 
+ WL_TK_ACT[490] WL_TK_ACT[491] WL_TK_ACT[492] WL_TK_ACT[493] WL_TK_ACT[494] 
+ WL_TK_ACT[495] WL_TK_ACT[496] WL_TK_ACT[497] WL_TK_ACT[498] WL_TK_ACT[499] 
+ WL_TK_ACT[500] WL_TK_ACT[501] WL_TK_ACT[502] WL_TK_ACT[503] WL_TK_ACT[504] 
+ WL_TK_ACT[505] WL_TK_ACT[506] WL_TK_ACT[507] WL_TK_ACT[508] WL_TK_ACT[509] 
+ WL_TK_ACT[510] WL_TK_ACT[511] WL_TK_LD WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] 
+ X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] 
+ XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YM[0] YM[1] YM[2] 
+ YM[3]
*.PININFO AWT:I BIST:I BWEBM_LL:I BWEBM_LR:I BWEB_LL:I BWEB_LR:I CEB:I CEBM:I 
*.PININFO CLK:I DM_LL:I DM_LR:I D_LL:I D_LR:I FAD1[0]:I FAD1[1]:I FAD1[2]:I 
*.PININFO FAD1[3]:I FAD1[4]:I FAD1[5]:I FAD1[6]:I FAD1[7]:I FAD1[8]:I 
*.PININFO FAD1[9]:I FAD1[10]:I FAD2[0]:I FAD2[1]:I FAD2[2]:I FAD2[3]:I 
*.PININFO FAD2[4]:I FAD2[5]:I FAD2[6]:I FAD2[7]:I FAD2[8]:I FAD2[9]:I 
*.PININFO FAD2[10]:I PD:I PTSEL:I REDEN1:I REDEN2:I RSTB:I RTSEL[0]:I 
*.PININFO RTSEL[1]:I SCLK:I SDIN:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I 
*.PININFO XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I 
*.PININFO Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I Q_LL:O Q_LR:O SDOUT:O 
*.PININFO VDDI:B VSSI:B WL_TK_ACT[0]:B WL_TK_ACT[1]:B WL_TK_ACT[2]:B 
*.PININFO WL_TK_ACT[3]:B WL_TK_ACT[4]:B WL_TK_ACT[5]:B WL_TK_ACT[6]:B 
*.PININFO WL_TK_ACT[7]:B WL_TK_ACT[8]:B WL_TK_ACT[9]:B WL_TK_ACT[10]:B 
*.PININFO WL_TK_ACT[11]:B WL_TK_ACT[12]:B WL_TK_ACT[13]:B WL_TK_ACT[14]:B 
*.PININFO WL_TK_ACT[15]:B WL_TK_ACT[16]:B WL_TK_ACT[17]:B WL_TK_ACT[18]:B 
*.PININFO WL_TK_ACT[19]:B WL_TK_ACT[20]:B WL_TK_ACT[21]:B WL_TK_ACT[22]:B 
*.PININFO WL_TK_ACT[23]:B WL_TK_ACT[24]:B WL_TK_ACT[25]:B WL_TK_ACT[26]:B 
*.PININFO WL_TK_ACT[27]:B WL_TK_ACT[28]:B WL_TK_ACT[29]:B WL_TK_ACT[30]:B 
*.PININFO WL_TK_ACT[31]:B WL_TK_ACT[32]:B WL_TK_ACT[33]:B WL_TK_ACT[34]:B 
*.PININFO WL_TK_ACT[35]:B WL_TK_ACT[36]:B WL_TK_ACT[37]:B WL_TK_ACT[38]:B 
*.PININFO WL_TK_ACT[39]:B WL_TK_ACT[40]:B WL_TK_ACT[41]:B WL_TK_ACT[42]:B 
*.PININFO WL_TK_ACT[43]:B WL_TK_ACT[44]:B WL_TK_ACT[45]:B WL_TK_ACT[46]:B 
*.PININFO WL_TK_ACT[47]:B WL_TK_ACT[48]:B WL_TK_ACT[49]:B WL_TK_ACT[50]:B 
*.PININFO WL_TK_ACT[51]:B WL_TK_ACT[52]:B WL_TK_ACT[53]:B WL_TK_ACT[54]:B 
*.PININFO WL_TK_ACT[55]:B WL_TK_ACT[56]:B WL_TK_ACT[57]:B WL_TK_ACT[58]:B 
*.PININFO WL_TK_ACT[59]:B WL_TK_ACT[60]:B WL_TK_ACT[61]:B WL_TK_ACT[62]:B 
*.PININFO WL_TK_ACT[63]:B WL_TK_ACT[64]:B WL_TK_ACT[65]:B WL_TK_ACT[66]:B 
*.PININFO WL_TK_ACT[67]:B WL_TK_ACT[68]:B WL_TK_ACT[69]:B WL_TK_ACT[70]:B 
*.PININFO WL_TK_ACT[71]:B WL_TK_ACT[72]:B WL_TK_ACT[73]:B WL_TK_ACT[74]:B 
*.PININFO WL_TK_ACT[75]:B WL_TK_ACT[76]:B WL_TK_ACT[77]:B WL_TK_ACT[78]:B 
*.PININFO WL_TK_ACT[79]:B WL_TK_ACT[80]:B WL_TK_ACT[81]:B WL_TK_ACT[82]:B 
*.PININFO WL_TK_ACT[83]:B WL_TK_ACT[84]:B WL_TK_ACT[85]:B WL_TK_ACT[86]:B 
*.PININFO WL_TK_ACT[87]:B WL_TK_ACT[88]:B WL_TK_ACT[89]:B WL_TK_ACT[90]:B 
*.PININFO WL_TK_ACT[91]:B WL_TK_ACT[92]:B WL_TK_ACT[93]:B WL_TK_ACT[94]:B 
*.PININFO WL_TK_ACT[95]:B WL_TK_ACT[96]:B WL_TK_ACT[97]:B WL_TK_ACT[98]:B 
*.PININFO WL_TK_ACT[99]:B WL_TK_ACT[100]:B WL_TK_ACT[101]:B WL_TK_ACT[102]:B 
*.PININFO WL_TK_ACT[103]:B WL_TK_ACT[104]:B WL_TK_ACT[105]:B WL_TK_ACT[106]:B 
*.PININFO WL_TK_ACT[107]:B WL_TK_ACT[108]:B WL_TK_ACT[109]:B WL_TK_ACT[110]:B 
*.PININFO WL_TK_ACT[111]:B WL_TK_ACT[112]:B WL_TK_ACT[113]:B WL_TK_ACT[114]:B 
*.PININFO WL_TK_ACT[115]:B WL_TK_ACT[116]:B WL_TK_ACT[117]:B WL_TK_ACT[118]:B 
*.PININFO WL_TK_ACT[119]:B WL_TK_ACT[120]:B WL_TK_ACT[121]:B WL_TK_ACT[122]:B 
*.PININFO WL_TK_ACT[123]:B WL_TK_ACT[124]:B WL_TK_ACT[125]:B WL_TK_ACT[126]:B 
*.PININFO WL_TK_ACT[127]:B WL_TK_ACT[128]:B WL_TK_ACT[129]:B WL_TK_ACT[130]:B 
*.PININFO WL_TK_ACT[131]:B WL_TK_ACT[132]:B WL_TK_ACT[133]:B WL_TK_ACT[134]:B 
*.PININFO WL_TK_ACT[135]:B WL_TK_ACT[136]:B WL_TK_ACT[137]:B WL_TK_ACT[138]:B 
*.PININFO WL_TK_ACT[139]:B WL_TK_ACT[140]:B WL_TK_ACT[141]:B WL_TK_ACT[142]:B 
*.PININFO WL_TK_ACT[143]:B WL_TK_ACT[144]:B WL_TK_ACT[145]:B WL_TK_ACT[146]:B 
*.PININFO WL_TK_ACT[147]:B WL_TK_ACT[148]:B WL_TK_ACT[149]:B WL_TK_ACT[150]:B 
*.PININFO WL_TK_ACT[151]:B WL_TK_ACT[152]:B WL_TK_ACT[153]:B WL_TK_ACT[154]:B 
*.PININFO WL_TK_ACT[155]:B WL_TK_ACT[156]:B WL_TK_ACT[157]:B WL_TK_ACT[158]:B 
*.PININFO WL_TK_ACT[159]:B WL_TK_ACT[160]:B WL_TK_ACT[161]:B WL_TK_ACT[162]:B 
*.PININFO WL_TK_ACT[163]:B WL_TK_ACT[164]:B WL_TK_ACT[165]:B WL_TK_ACT[166]:B 
*.PININFO WL_TK_ACT[167]:B WL_TK_ACT[168]:B WL_TK_ACT[169]:B WL_TK_ACT[170]:B 
*.PININFO WL_TK_ACT[171]:B WL_TK_ACT[172]:B WL_TK_ACT[173]:B WL_TK_ACT[174]:B 
*.PININFO WL_TK_ACT[175]:B WL_TK_ACT[176]:B WL_TK_ACT[177]:B WL_TK_ACT[178]:B 
*.PININFO WL_TK_ACT[179]:B WL_TK_ACT[180]:B WL_TK_ACT[181]:B WL_TK_ACT[182]:B 
*.PININFO WL_TK_ACT[183]:B WL_TK_ACT[184]:B WL_TK_ACT[185]:B WL_TK_ACT[186]:B 
*.PININFO WL_TK_ACT[187]:B WL_TK_ACT[188]:B WL_TK_ACT[189]:B WL_TK_ACT[190]:B 
*.PININFO WL_TK_ACT[191]:B WL_TK_ACT[192]:B WL_TK_ACT[193]:B WL_TK_ACT[194]:B 
*.PININFO WL_TK_ACT[195]:B WL_TK_ACT[196]:B WL_TK_ACT[197]:B WL_TK_ACT[198]:B 
*.PININFO WL_TK_ACT[199]:B WL_TK_ACT[200]:B WL_TK_ACT[201]:B WL_TK_ACT[202]:B 
*.PININFO WL_TK_ACT[203]:B WL_TK_ACT[204]:B WL_TK_ACT[205]:B WL_TK_ACT[206]:B 
*.PININFO WL_TK_ACT[207]:B WL_TK_ACT[208]:B WL_TK_ACT[209]:B WL_TK_ACT[210]:B 
*.PININFO WL_TK_ACT[211]:B WL_TK_ACT[212]:B WL_TK_ACT[213]:B WL_TK_ACT[214]:B 
*.PININFO WL_TK_ACT[215]:B WL_TK_ACT[216]:B WL_TK_ACT[217]:B WL_TK_ACT[218]:B 
*.PININFO WL_TK_ACT[219]:B WL_TK_ACT[220]:B WL_TK_ACT[221]:B WL_TK_ACT[222]:B 
*.PININFO WL_TK_ACT[223]:B WL_TK_ACT[224]:B WL_TK_ACT[225]:B WL_TK_ACT[226]:B 
*.PININFO WL_TK_ACT[227]:B WL_TK_ACT[228]:B WL_TK_ACT[229]:B WL_TK_ACT[230]:B 
*.PININFO WL_TK_ACT[231]:B WL_TK_ACT[232]:B WL_TK_ACT[233]:B WL_TK_ACT[234]:B 
*.PININFO WL_TK_ACT[235]:B WL_TK_ACT[236]:B WL_TK_ACT[237]:B WL_TK_ACT[238]:B 
*.PININFO WL_TK_ACT[239]:B WL_TK_ACT[240]:B WL_TK_ACT[241]:B WL_TK_ACT[242]:B 
*.PININFO WL_TK_ACT[243]:B WL_TK_ACT[244]:B WL_TK_ACT[245]:B WL_TK_ACT[246]:B 
*.PININFO WL_TK_ACT[247]:B WL_TK_ACT[248]:B WL_TK_ACT[249]:B WL_TK_ACT[250]:B 
*.PININFO WL_TK_ACT[251]:B WL_TK_ACT[252]:B WL_TK_ACT[253]:B WL_TK_ACT[254]:B 
*.PININFO WL_TK_ACT[255]:B WL_TK_ACT[256]:B WL_TK_ACT[257]:B WL_TK_ACT[258]:B 
*.PININFO WL_TK_ACT[259]:B WL_TK_ACT[260]:B WL_TK_ACT[261]:B WL_TK_ACT[262]:B 
*.PININFO WL_TK_ACT[263]:B WL_TK_ACT[264]:B WL_TK_ACT[265]:B WL_TK_ACT[266]:B 
*.PININFO WL_TK_ACT[267]:B WL_TK_ACT[268]:B WL_TK_ACT[269]:B WL_TK_ACT[270]:B 
*.PININFO WL_TK_ACT[271]:B WL_TK_ACT[272]:B WL_TK_ACT[273]:B WL_TK_ACT[274]:B 
*.PININFO WL_TK_ACT[275]:B WL_TK_ACT[276]:B WL_TK_ACT[277]:B WL_TK_ACT[278]:B 
*.PININFO WL_TK_ACT[279]:B WL_TK_ACT[280]:B WL_TK_ACT[281]:B WL_TK_ACT[282]:B 
*.PININFO WL_TK_ACT[283]:B WL_TK_ACT[284]:B WL_TK_ACT[285]:B WL_TK_ACT[286]:B 
*.PININFO WL_TK_ACT[287]:B WL_TK_ACT[288]:B WL_TK_ACT[289]:B WL_TK_ACT[290]:B 
*.PININFO WL_TK_ACT[291]:B WL_TK_ACT[292]:B WL_TK_ACT[293]:B WL_TK_ACT[294]:B 
*.PININFO WL_TK_ACT[295]:B WL_TK_ACT[296]:B WL_TK_ACT[297]:B WL_TK_ACT[298]:B 
*.PININFO WL_TK_ACT[299]:B WL_TK_ACT[300]:B WL_TK_ACT[301]:B WL_TK_ACT[302]:B 
*.PININFO WL_TK_ACT[303]:B WL_TK_ACT[304]:B WL_TK_ACT[305]:B WL_TK_ACT[306]:B 
*.PININFO WL_TK_ACT[307]:B WL_TK_ACT[308]:B WL_TK_ACT[309]:B WL_TK_ACT[310]:B 
*.PININFO WL_TK_ACT[311]:B WL_TK_ACT[312]:B WL_TK_ACT[313]:B WL_TK_ACT[314]:B 
*.PININFO WL_TK_ACT[315]:B WL_TK_ACT[316]:B WL_TK_ACT[317]:B WL_TK_ACT[318]:B 
*.PININFO WL_TK_ACT[319]:B WL_TK_ACT[320]:B WL_TK_ACT[321]:B WL_TK_ACT[322]:B 
*.PININFO WL_TK_ACT[323]:B WL_TK_ACT[324]:B WL_TK_ACT[325]:B WL_TK_ACT[326]:B 
*.PININFO WL_TK_ACT[327]:B WL_TK_ACT[328]:B WL_TK_ACT[329]:B WL_TK_ACT[330]:B 
*.PININFO WL_TK_ACT[331]:B WL_TK_ACT[332]:B WL_TK_ACT[333]:B WL_TK_ACT[334]:B 
*.PININFO WL_TK_ACT[335]:B WL_TK_ACT[336]:B WL_TK_ACT[337]:B WL_TK_ACT[338]:B 
*.PININFO WL_TK_ACT[339]:B WL_TK_ACT[340]:B WL_TK_ACT[341]:B WL_TK_ACT[342]:B 
*.PININFO WL_TK_ACT[343]:B WL_TK_ACT[344]:B WL_TK_ACT[345]:B WL_TK_ACT[346]:B 
*.PININFO WL_TK_ACT[347]:B WL_TK_ACT[348]:B WL_TK_ACT[349]:B WL_TK_ACT[350]:B 
*.PININFO WL_TK_ACT[351]:B WL_TK_ACT[352]:B WL_TK_ACT[353]:B WL_TK_ACT[354]:B 
*.PININFO WL_TK_ACT[355]:B WL_TK_ACT[356]:B WL_TK_ACT[357]:B WL_TK_ACT[358]:B 
*.PININFO WL_TK_ACT[359]:B WL_TK_ACT[360]:B WL_TK_ACT[361]:B WL_TK_ACT[362]:B 
*.PININFO WL_TK_ACT[363]:B WL_TK_ACT[364]:B WL_TK_ACT[365]:B WL_TK_ACT[366]:B 
*.PININFO WL_TK_ACT[367]:B WL_TK_ACT[368]:B WL_TK_ACT[369]:B WL_TK_ACT[370]:B 
*.PININFO WL_TK_ACT[371]:B WL_TK_ACT[372]:B WL_TK_ACT[373]:B WL_TK_ACT[374]:B 
*.PININFO WL_TK_ACT[375]:B WL_TK_ACT[376]:B WL_TK_ACT[377]:B WL_TK_ACT[378]:B 
*.PININFO WL_TK_ACT[379]:B WL_TK_ACT[380]:B WL_TK_ACT[381]:B WL_TK_ACT[382]:B 
*.PININFO WL_TK_ACT[383]:B WL_TK_ACT[384]:B WL_TK_ACT[385]:B WL_TK_ACT[386]:B 
*.PININFO WL_TK_ACT[387]:B WL_TK_ACT[388]:B WL_TK_ACT[389]:B WL_TK_ACT[390]:B 
*.PININFO WL_TK_ACT[391]:B WL_TK_ACT[392]:B WL_TK_ACT[393]:B WL_TK_ACT[394]:B 
*.PININFO WL_TK_ACT[395]:B WL_TK_ACT[396]:B WL_TK_ACT[397]:B WL_TK_ACT[398]:B 
*.PININFO WL_TK_ACT[399]:B WL_TK_ACT[400]:B WL_TK_ACT[401]:B WL_TK_ACT[402]:B 
*.PININFO WL_TK_ACT[403]:B WL_TK_ACT[404]:B WL_TK_ACT[405]:B WL_TK_ACT[406]:B 
*.PININFO WL_TK_ACT[407]:B WL_TK_ACT[408]:B WL_TK_ACT[409]:B WL_TK_ACT[410]:B 
*.PININFO WL_TK_ACT[411]:B WL_TK_ACT[412]:B WL_TK_ACT[413]:B WL_TK_ACT[414]:B 
*.PININFO WL_TK_ACT[415]:B WL_TK_ACT[416]:B WL_TK_ACT[417]:B WL_TK_ACT[418]:B 
*.PININFO WL_TK_ACT[419]:B WL_TK_ACT[420]:B WL_TK_ACT[421]:B WL_TK_ACT[422]:B 
*.PININFO WL_TK_ACT[423]:B WL_TK_ACT[424]:B WL_TK_ACT[425]:B WL_TK_ACT[426]:B 
*.PININFO WL_TK_ACT[427]:B WL_TK_ACT[428]:B WL_TK_ACT[429]:B WL_TK_ACT[430]:B 
*.PININFO WL_TK_ACT[431]:B WL_TK_ACT[432]:B WL_TK_ACT[433]:B WL_TK_ACT[434]:B 
*.PININFO WL_TK_ACT[435]:B WL_TK_ACT[436]:B WL_TK_ACT[437]:B WL_TK_ACT[438]:B 
*.PININFO WL_TK_ACT[439]:B WL_TK_ACT[440]:B WL_TK_ACT[441]:B WL_TK_ACT[442]:B 
*.PININFO WL_TK_ACT[443]:B WL_TK_ACT[444]:B WL_TK_ACT[445]:B WL_TK_ACT[446]:B 
*.PININFO WL_TK_ACT[447]:B WL_TK_ACT[448]:B WL_TK_ACT[449]:B WL_TK_ACT[450]:B 
*.PININFO WL_TK_ACT[451]:B WL_TK_ACT[452]:B WL_TK_ACT[453]:B WL_TK_ACT[454]:B 
*.PININFO WL_TK_ACT[455]:B WL_TK_ACT[456]:B WL_TK_ACT[457]:B WL_TK_ACT[458]:B 
*.PININFO WL_TK_ACT[459]:B WL_TK_ACT[460]:B WL_TK_ACT[461]:B WL_TK_ACT[462]:B 
*.PININFO WL_TK_ACT[463]:B WL_TK_ACT[464]:B WL_TK_ACT[465]:B WL_TK_ACT[466]:B 
*.PININFO WL_TK_ACT[467]:B WL_TK_ACT[468]:B WL_TK_ACT[469]:B WL_TK_ACT[470]:B 
*.PININFO WL_TK_ACT[471]:B WL_TK_ACT[472]:B WL_TK_ACT[473]:B WL_TK_ACT[474]:B 
*.PININFO WL_TK_ACT[475]:B WL_TK_ACT[476]:B WL_TK_ACT[477]:B WL_TK_ACT[478]:B 
*.PININFO WL_TK_ACT[479]:B WL_TK_ACT[480]:B WL_TK_ACT[481]:B WL_TK_ACT[482]:B 
*.PININFO WL_TK_ACT[483]:B WL_TK_ACT[484]:B WL_TK_ACT[485]:B WL_TK_ACT[486]:B 
*.PININFO WL_TK_ACT[487]:B WL_TK_ACT[488]:B WL_TK_ACT[489]:B WL_TK_ACT[490]:B 
*.PININFO WL_TK_ACT[491]:B WL_TK_ACT[492]:B WL_TK_ACT[493]:B WL_TK_ACT[494]:B 
*.PININFO WL_TK_ACT[495]:B WL_TK_ACT[496]:B WL_TK_ACT[497]:B WL_TK_ACT[498]:B 
*.PININFO WL_TK_ACT[499]:B WL_TK_ACT[500]:B WL_TK_ACT[501]:B WL_TK_ACT[502]:B 
*.PININFO WL_TK_ACT[503]:B WL_TK_ACT[504]:B WL_TK_ACT[505]:B WL_TK_ACT[506]:B 
*.PININFO WL_TK_ACT[507]:B WL_TK_ACT[508]:B WL_TK_ACT[509]:B WL_TK_ACT[510]:B 
*.PININFO WL_TK_ACT[511]:B WL_TK_LD:B
XBK_WLDV_U VDDHD VDDI DEC_X0_7[0] DEC_X0_7[1] DEC_X0_7[2] DEC_X0_7[3] 
+ DEC_X0_7[4] DEC_X0_7[5] DEC_X0_7[6] DEC_X0_7[7] NET0103[0] NET0103[1] 
+ NET0103[2] NET0103[3] NET0103[4] NET0103[5] NET0103[6] NET0103[7] 
+ DEC_X1_7[0] DEC_X1_7[1] DEC_X1_7[2] DEC_X1_7[3] DEC_X1_7[4] DEC_X1_7[5] 
+ DEC_X1_7[6] DEC_X1_7[7] NET0102[0] NET0102[1] NET0102[2] NET0102[3] 
+ NET0102[4] NET0102[5] NET0102[6] NET0102[7] DEC_X2_7[0] DEC_X2_7[1] 
+ DEC_X2_7[2] DEC_X2_7[3] NET097[0] NET097[1] NET097[2] NET097[3] DEC_X3_7[0] 
+ DEC_X3_7[1] DEC_X3_7[2] DEC_X3_7[3] DEC_X3_7[4] DEC_X3_7[5] DEC_X3_7[6] 
+ DEC_X3_7[7] NET0100[0] NET0100[1] NET0100[2] NET0100[3] NET0100[4] 
+ NET0100[5] NET0100[6] NET0100[7] DEC_Y_7[0] DEC_Y_7[1] DEC_Y_7[2] DEC_Y_7[3] 
+ DEC_Y_7[4] DEC_Y_7[5] DEC_Y_7[6] DEC_Y_7[7] NET0121[0] NET0121[1] NET0121[2] 
+ NET0121[3] NET0121[4] NET0121[5] NET0121[6] NET0121[7] PD_BUF_7 NET0107 
+ PD_CVDDBUF_7 NET0106 RW_RE_7 NET0105 VDDHD VDDI VSSI WLPYB_7 NET897 WLPY_7 
+ NET915 WLP_SAE_7 WLP_SAE_TK_7 WLP_SAE_TK_8 WLP_SAE_8 WL_LU1[0] WL_LU1[1] 
+ WL_RU1[0] WL_RU1[1] YL_7[0] NET0111 S1AHSF400W40_BK_WLDV_U_SIM
XBK_WLDV_D VDDHD VDDI DEC_X0_1[0] DEC_X0_1[1] DEC_X0_1[2] DEC_X0_1[3] 
+ DEC_X0_1[4] DEC_X0_1[5] DEC_X0_1[6] DEC_X0_1[7] DEC_X0_2[0] DEC_X0_2[1] 
+ DEC_X0_2[2] DEC_X0_2[3] DEC_X0_2[4] DEC_X0_2[5] DEC_X0_2[6] DEC_X0_2[7] 
+ DEC_X1_1[0] DEC_X1_1[1] DEC_X1_1[2] DEC_X1_1[3] DEC_X1_1[4] DEC_X1_1[5] 
+ DEC_X1_1[6] DEC_X1_1[7] DEC_X1_2[0] DEC_X1_2[1] DEC_X1_2[2] DEC_X1_2[3] 
+ DEC_X1_2[4] DEC_X1_2[5] DEC_X1_2[6] DEC_X1_2[7] DEC_X2_1[0] DEC_X2_1[1] 
+ DEC_X2_1[2] DEC_X2_1[3] DEC_X2_2[0] DEC_X2_2[1] DEC_X2_2[2] DEC_X2_2[3] 
+ DEC_X3_1[0] DEC_X3_1[1] DEC_X3_1[2] DEC_X3_1[3] DEC_X3_1[4] DEC_X3_1[5] 
+ DEC_X3_1[6] DEC_X3_1[7] DEC_X3_2[0] DEC_X3_2[1] DEC_X3_2[2] DEC_X3_2[3] 
+ DEC_X3_2[4] DEC_X3_2[5] DEC_X3_2[6] DEC_X3_2[7] DEC_Y_1[0] DEC_Y_1[1] 
+ DEC_Y_1[2] DEC_Y_1[3] DEC_Y_1[4] DEC_Y_1[5] DEC_Y_1[6] DEC_Y_1[7] DEC_Y_2[0] 
+ DEC_Y_2[1] DEC_Y_2[2] DEC_Y_2[3] DEC_Y_2[4] DEC_Y_2[5] DEC_Y_2[6] DEC_Y_2[7] 
+ PD_BUF_1 PD_BUF_2 PD_CVDDBUF_1 PD_CVDDBUF_2 RW_RE_1 RW_RE_2 VDDHD VDDI VSSI 
+ NET124 WLPYB_2 NET125 WLPY_2 WLP_SAE_1 WLP_SAE_TK_1 WLP_SAE_TK_2 WLP_SAE_2 
+ WL_LD1[0] WL_LD1[1] WL_RD1[0] WL_RD1[1] YL_1[0] YL_2[0] S1AHSF400W40_BK_WLDV_D_SIM
XWLPY_LD_U VDDHD VDDI VDDHD VDDI VSSI WLPYB_4 WLPYB_7 WLPY_4 WLPY_7 
+ S1AHSF400W40_WLPY_LD_SIM
XWLPY_LD_D VDDHD VDDI VDDHD VDDI VSSI WLPYB_2 WLPYB_3 WLPY_2 WLPY_3 
+ S1AHSF400W40_WLPY_LD_SIM
XBK_LCNT_D BLEQ_DN_LD1 BLEQ_DN_RD1 BLEQ_UP_LD1 BLEQ_UP_RD1 VDDHD VDDI 
+ DEC_X0_3[0] DEC_X0_3[1] DEC_X0_3[2] DEC_X0_3[3] DEC_X0_3[4] DEC_X0_3[5] 
+ DEC_X0_3[6] DEC_X0_3[7] DEC_X0_4[0] DEC_X0_4[1] DEC_X0_4[2] DEC_X0_4[3] 
+ DEC_X0_4[4] DEC_X0_4[5] DEC_X0_4[6] DEC_X0_4[7] DEC_X1_3[0] DEC_X1_3[1] 
+ DEC_X1_3[2] DEC_X1_3[3] DEC_X1_3[4] DEC_X1_3[5] DEC_X1_3[6] DEC_X1_3[7] 
+ DEC_X1_4[0] DEC_X1_4[1] DEC_X1_4[2] DEC_X1_4[3] DEC_X1_4[4] DEC_X1_4[5] 
+ DEC_X1_4[6] DEC_X1_4[7] DEC_X2_3[0] DEC_X2_3[1] DEC_X2_3[2] DEC_X2_3[3] 
+ DEC_X2_4[0] DEC_X2_4[1] DEC_X2_4[2] DEC_X2_4[3] DEC_X3_3[0] DEC_X3_3[1] 
+ DEC_X3_3[2] DEC_X3_3[3] DEC_X3_3[4] DEC_X3_3[5] DEC_X3_3[6] DEC_X3_3[7] 
+ DEC_X3_4[0] DEC_X3_4[1] DEC_X3_4[2] DEC_X3_4[3] DEC_X3_4[4] DEC_X3_4[5] 
+ DEC_X3_4[6] DEC_X3_4[7] DEC_Y_3[0] DEC_Y_3[1] DEC_Y_3[2] DEC_Y_3[3] 
+ DEC_Y_3[4] DEC_Y_3[5] DEC_Y_3[6] DEC_Y_3[7] Y_DN_LD1[0] Y_DN_LD1[1] 
+ Y_DN_LD1[2] Y_DN_LD1[3] Y_DN_LD1[4] Y_DN_LD1[5] Y_DN_LD1[6] Y_DN_LD1[7] 
+ Y_DN_RD1[0] Y_DN_RD1[1] Y_DN_RD1[2] Y_DN_RD1[3] Y_DN_RD1[4] Y_DN_RD1[5] 
+ Y_DN_RD1[6] Y_DN_RD1[7] DEC_Y_4[0] DEC_Y_4[1] DEC_Y_4[2] DEC_Y_4[3] 
+ DEC_Y_4[4] DEC_Y_4[5] DEC_Y_4[6] DEC_Y_4[7] Y_UP_LD1[0] Y_UP_LD1[1] 
+ Y_UP_LD1[2] Y_UP_LD1[3] Y_UP_LD1[4] Y_UP_LD1[5] Y_UP_LD1[6] Y_UP_LD1[7] 
+ Y_UP_RD1[0] Y_UP_RD1[1] Y_UP_RD1[2] Y_UP_RD1[3] Y_UP_RD1[4] Y_UP_RD1[5] 
+ Y_UP_RD1[6] Y_UP_RD1[7] PD_BUF_3 PD_BUF_4 PD_CVDDBUF_3 PD_CVDDBUF_4 RE_LD1 
+ RE_RD1 RW_RE_3 RW_RE_4 SAEB_LD1 SAEB_RD1 VDDHD VDDI VSSI WE_LD1 WE_RD1 
+ WLPYB_3 WLPYB_4 WLPY_3 WLPY_4 WLP_SAE_3 WLP_SAE_TK_3 WLP_SAE_TK_4 WLP_SAE_4 
+ YL_3[0] YL_LD1[0] YL_LD1[1] YL_RD1[0] YL_RD1[1] YL_4[0] S1AHSF400W40_BK_LCNT_D_SIM
XBK_WLDV_LD_D VDDHD VDDI DEC_X0_2[0] DEC_X0_2[1] DEC_X0_2[2] DEC_X0_2[3] 
+ DEC_X0_2[4] DEC_X0_2[5] DEC_X0_2[6] DEC_X0_2[7] DEC_X0_3[0] DEC_X0_3[1] 
+ DEC_X0_3[2] DEC_X0_3[3] DEC_X0_3[4] DEC_X0_3[5] DEC_X0_3[6] DEC_X0_3[7] 
+ DEC_X1_2[0] DEC_X1_2[1] DEC_X1_2[2] DEC_X1_2[3] DEC_X1_2[4] DEC_X1_2[5] 
+ DEC_X1_2[6] DEC_X1_2[7] DEC_X1_3[0] DEC_X1_3[1] DEC_X1_3[2] DEC_X1_3[3] 
+ DEC_X1_3[4] DEC_X1_3[5] DEC_X1_3[6] DEC_X1_3[7] DEC_X2_2[0] DEC_X2_2[1] 
+ DEC_X2_2[2] DEC_X2_2[3] DEC_X2_3[0] DEC_X2_3[1] DEC_X2_3[2] DEC_X2_3[3] 
+ DEC_X3_2[0] DEC_X3_2[1] DEC_X3_2[2] DEC_X3_2[3] DEC_X3_2[4] DEC_X3_2[5] 
+ DEC_X3_2[6] DEC_X3_2[7] DEC_X3_3[0] DEC_X3_3[1] DEC_X3_3[2] DEC_X3_3[3] 
+ DEC_X3_3[4] DEC_X3_3[5] DEC_X3_3[6] DEC_X3_3[7] DEC_Y_2[0] DEC_Y_2[1] 
+ DEC_Y_2[2] DEC_Y_2[3] DEC_Y_2[4] DEC_Y_2[5] DEC_Y_2[6] DEC_Y_2[7] DEC_Y_3[0] 
+ DEC_Y_3[1] DEC_Y_3[2] DEC_Y_3[3] DEC_Y_3[4] DEC_Y_3[5] DEC_Y_3[6] DEC_Y_3[7] 
+ PD_BUF_2 PD_BUF_3 PD_CVDDBUF_2 PD_CVDDBUF_3 RW_RE_2 RW_RE_3 VDDHD VDDI VSSI 
+ WLP_SAE_2 WLP_SAE_TK_2 WLP_SAE_TK_3 WLP_SAE_3 YL_2[0] YL_3[0] 
+ S1AHSF400W40_BK_WLDV_LD_SIM
XBK_WLDV_LD_U VDDHD VDDI DEC_X0_4[0] DEC_X0_4[1] DEC_X0_4[2] DEC_X0_4[3] 
+ DEC_X0_4[4] DEC_X0_4[5] DEC_X0_4[6] DEC_X0_4[7] DEC_X0_7[0] DEC_X0_7[1] 
+ DEC_X0_7[2] DEC_X0_7[3] DEC_X0_7[4] DEC_X0_7[5] DEC_X0_7[6] DEC_X0_7[7] 
+ DEC_X1_4[0] DEC_X1_4[1] DEC_X1_4[2] DEC_X1_4[3] DEC_X1_4[4] DEC_X1_4[5] 
+ DEC_X1_4[6] DEC_X1_4[7] DEC_X1_7[0] DEC_X1_7[1] DEC_X1_7[2] DEC_X1_7[3] 
+ DEC_X1_7[4] DEC_X1_7[5] DEC_X1_7[6] DEC_X1_7[7] DEC_X2_4[0] DEC_X2_4[1] 
+ DEC_X2_4[2] DEC_X2_4[3] DEC_X2_7[0] DEC_X2_7[1] DEC_X2_7[2] DEC_X2_7[3] 
+ DEC_X3_4[0] DEC_X3_4[1] DEC_X3_4[2] DEC_X3_4[3] DEC_X3_4[4] DEC_X3_4[5] 
+ DEC_X3_4[6] DEC_X3_4[7] DEC_X3_7[0] DEC_X3_7[1] DEC_X3_7[2] DEC_X3_7[3] 
+ DEC_X3_7[4] DEC_X3_7[5] DEC_X3_7[6] DEC_X3_7[7] DEC_Y_4[0] DEC_Y_4[1] 
+ DEC_Y_4[2] DEC_Y_4[3] DEC_Y_4[4] DEC_Y_4[5] DEC_Y_4[6] DEC_Y_4[7] DEC_Y_7[0] 
+ DEC_Y_7[1] DEC_Y_7[2] DEC_Y_7[3] DEC_Y_7[4] DEC_Y_7[5] DEC_Y_7[6] DEC_Y_7[7] 
+ PD_BUF_4 PD_BUF_7 PD_CVDDBUF_4 PD_CVDDBUF_7 RW_RE_4 RW_RE_7 VDDHD VDDI VSSI 
+ WLP_SAE_4 WLP_SAE_TK_4 WLP_SAE_TK_7 WLP_SAE_7 YL_4[0] YL_7[0] 
+ S1AHSF400W40_BK_WLDV_LD_SIM
XTRKPRE PD TRKBL WL_TK VDDHD VDDI VSSI TIEH_BT TIEL S1AHSF400W40_TRKPRE_SIM
XBK_TOP_EDGE VDDHD VDDI VSSI WLP_SAE_8 WLP_SAE_TK_8 S1AHSF400W40_BK_TOP_EDGE_SIM
XARR_LIO_LD_LD BLEQ_DN_LD3 BLEQ_DN_LD2 BLEQ_UP_LD3 BLEQ_UP_LD2 VDDI RE_LD3 
+ RE_LD2 SAEB_LD3 SAEB_LD2 VDDHD VDDI VSSI WE_LD3 WE_LD2 YL_LD3[0] YL_LD3[1] 
+ YL_LD2[0] YL_LD2[1] Y_DN_LD3[0] Y_DN_LD3[1] Y_DN_LD3[2] Y_DN_LD3[3] 
+ Y_DN_LD3[4] Y_DN_LD3[5] Y_DN_LD3[6] Y_DN_LD3[7] Y_DN_LD2[0] Y_DN_LD2[1] 
+ Y_DN_LD2[2] Y_DN_LD2[3] Y_DN_LD2[4] Y_DN_LD2[5] Y_DN_LD2[6] Y_DN_LD2[7] 
+ Y_UP_LD3[0] Y_UP_LD3[1] Y_UP_LD3[2] Y_UP_LD3[3] Y_UP_LD3[4] Y_UP_LD3[5] 
+ Y_UP_LD3[6] Y_UP_LD3[7] Y_UP_LD2[0] Y_UP_LD2[1] Y_UP_LD2[2] Y_UP_LD2[3] 
+ Y_UP_LD2[4] Y_UP_LD2[5] Y_UP_LD2[6] Y_UP_LD2[7] S1AHSF400W40_ARR_LIO_LD_SIM
XARR_LIO_LD_RD BLEQ_DN_RD2 BLEQ_DN_RD3 BLEQ_UP_RD2 BLEQ_UP_RD3 VDDI RE_RD2 
+ RE_RD3 SAEB_RD2 SAEB_RD3 VDDHD VDDI VSSI WE_RD2 WE_RD3 YL_RD2[0] YL_RD2[1] 
+ YL_RD3[0] YL_RD3[1] Y_DN_RD2[0] Y_DN_RD2[1] Y_DN_RD2[2] Y_DN_RD2[3] 
+ Y_DN_RD2[4] Y_DN_RD2[5] Y_DN_RD2[6] Y_DN_RD2[7] Y_DN_RD3[0] Y_DN_RD3[1] 
+ Y_DN_RD3[2] Y_DN_RD3[3] Y_DN_RD3[4] Y_DN_RD3[5] Y_DN_RD3[6] Y_DN_RD3[7] 
+ Y_UP_RD2[0] Y_UP_RD2[1] Y_UP_RD2[2] Y_UP_RD2[3] Y_UP_RD2[4] Y_UP_RD2[5] 
+ Y_UP_RD2[6] Y_UP_RD2[7] Y_UP_RD3[0] Y_UP_RD3[1] Y_UP_RD3[2] Y_UP_RD3[3] 
+ Y_UP_RD3[4] Y_UP_RD3[5] Y_UP_RD3[6] Y_UP_RD3[7] S1AHSF400W40_ARR_LIO_LD_SIM
XARR_LIO_LDR BLB_LR_3 BLB_DUM_LR_3 NET0324[0] NET0324[1] NET0324[2] NET0324[3] 
+ NET0324[4] NET0324[5] NET0324[6] NET0324[7] NET0324[8] NET0324[9] 
+ NET0324[10] NET0324[11] NET0324[12] NET0324[13] BLB_LR_4 BLB_DUM_LR_4 
+ NET0326[0] NET0326[1] NET0326[2] NET0326[3] NET0326[4] NET0326[5] NET0326[6] 
+ NET0326[7] NET0326[8] NET0326[9] NET0326[10] NET0326[11] NET0326[12] 
+ NET0326[13] BLEQ_DN_LD2 BLEQ_DN_LD1 BLEQ_UP_LD2 BLEQ_UP_LD1 BL_LR_3 
+ BL_DUM_LR_3 NET0329[0] NET0329[1] NET0329[2] NET0329[3] NET0329[4] 
+ NET0329[5] NET0329[6] NET0329[7] NET0329[8] NET0329[9] NET0329[10] 
+ NET0329[11] NET0329[12] NET0329[13] BL_LR_4 BL_DUM_LR_4 NET0327[0] 
+ NET0327[1] NET0327[2] NET0327[3] NET0327[4] NET0327[5] NET0327[6] NET0327[7] 
+ NET0327[8] NET0327[9] NET0327[10] NET0327[11] NET0327[12] NET0327[13] VDDI 
+ GBLB_LR_3 GBLB_LR_4 GBL_LR_3 GBL_LR_4 GWB_LR_3 GWB_LR_4 GW_LR_3 GW_LR_4 
+ RE_LD2 RE_LD1 SAEB_LD2 SAEB_LD1 VDDHD VDDI VSSI WE_LD2 WE_LD1 YL_LD2[0] 
+ YL_LD2[1] YL_LD1[0] YL_LD1[1] Y_DN_LD2[0] Y_DN_LD2[1] Y_DN_LD2[2] 
+ Y_DN_LD2[3] Y_DN_LD2[4] Y_DN_LD2[5] Y_DN_LD2[6] Y_DN_LD2[7] Y_DN_LD1[0] 
+ Y_DN_LD1[1] Y_DN_LD1[2] Y_DN_LD1[3] Y_DN_LD1[4] Y_DN_LD1[5] Y_DN_LD1[6] 
+ Y_DN_LD1[7] Y_UP_LD2[0] Y_UP_LD2[1] Y_UP_LD2[2] Y_UP_LD2[3] Y_UP_LD2[4] 
+ Y_UP_LD2[5] Y_UP_LD2[6] Y_UP_LD2[7] Y_UP_LD1[0] Y_UP_LD1[1] Y_UP_LD1[2] 
+ Y_UP_LD1[3] Y_UP_LD1[4] Y_UP_LD1[5] Y_UP_LD1[6] Y_UP_LD1[7] S1AHSF400W40_ARR_LIO_SIM
XARR_LIO_RDR NET363 NET0363 NET0364[0] NET0364[1] NET0364[2] NET0364[3] 
+ NET0364[4] NET0364[5] NET0364[6] NET0364[7] NET0364[8] NET0364[9] 
+ NET0364[10] NET0364[11] NET0364[12] NET0364[13] NET372 NET0365 NET0366[0] 
+ NET0366[1] NET0366[2] NET0366[3] NET0366[4] NET0366[5] NET0366[6] NET0366[7] 
+ NET0366[8] NET0366[9] NET0366[10] NET0366[11] NET0366[12] NET0366[13] 
+ BLEQ_DN_RD3 BLEQ_DN_RD4 BLEQ_UP_RD3 BLEQ_UP_RD4 NET371 NET0370 NET0369[0] 
+ NET0369[1] NET0369[2] NET0369[3] NET0369[4] NET0369[5] NET0369[6] NET0369[7] 
+ NET0369[8] NET0369[9] NET0369[10] NET0369[11] NET0369[12] NET0369[13] NET367 
+ NET0368 NET0367[0] NET0367[1] NET0367[2] NET0367[3] NET0367[4] NET0367[5] 
+ NET0367[6] NET0367[7] NET0367[8] NET0367[9] NET0367[10] NET0367[11] 
+ NET0367[12] NET0367[13] VDDI NET378 NET377 NET376 NET375 NET374 NET373 
+ NET370 NET369 RE_RD3 RE_RD4 SAEB_RD3 SAEB_RD4 VDDHD VDDI VSSI WE_RD3 WE_RD4 
+ YL_RD3[0] YL_RD3[1] YL_RD4[0] YL_RD4[1] Y_DN_RD3[0] Y_DN_RD3[1] Y_DN_RD3[2] 
+ Y_DN_RD3[3] Y_DN_RD3[4] Y_DN_RD3[5] Y_DN_RD3[6] Y_DN_RD3[7] Y_DN_RD4[0] 
+ Y_DN_RD4[1] Y_DN_RD4[2] Y_DN_RD4[3] Y_DN_RD4[4] Y_DN_RD4[5] Y_DN_RD4[6] 
+ Y_DN_RD4[7] Y_UP_RD3[0] Y_UP_RD3[1] Y_UP_RD3[2] Y_UP_RD3[3] Y_UP_RD3[4] 
+ Y_UP_RD3[5] Y_UP_RD3[6] Y_UP_RD3[7] Y_UP_RD4[0] Y_UP_RD4[1] Y_UP_RD4[2] 
+ Y_UP_RD4[3] Y_UP_RD4[4] Y_UP_RD4[5] Y_UP_RD4[6] Y_UP_RD4[7] S1AHSF400W40_ARR_LIO_SIM
XARR_LIO_RDL NET888 NET0403 NET0404[0] NET0404[1] NET0404[2] NET0404[3] 
+ NET0404[4] NET0404[5] NET0404[6] NET0404[7] NET0404[8] NET0404[9] 
+ NET0404[10] NET0404[11] NET0404[12] NET0404[13] NET868 NET0405 NET0406[0] 
+ NET0406[1] NET0406[2] NET0406[3] NET0406[4] NET0406[5] NET0406[6] NET0406[7] 
+ NET0406[8] NET0406[9] NET0406[10] NET0406[11] NET0406[12] NET0406[13] 
+ BLEQ_DN_RD1 BLEQ_DN_RD2 BLEQ_UP_RD1 BLEQ_UP_RD2 NET938 NET0410 NET0409[0] 
+ NET0409[1] NET0409[2] NET0409[3] NET0409[4] NET0409[5] NET0409[6] NET0409[7] 
+ NET0409[8] NET0409[9] NET0409[10] NET0409[11] NET0409[12] NET0409[13] NET883 
+ NET0408 NET0407[0] NET0407[1] NET0407[2] NET0407[3] NET0407[4] NET0407[5] 
+ NET0407[6] NET0407[7] NET0407[8] NET0407[9] NET0407[10] NET0407[11] 
+ NET0407[12] NET0407[13] VDDI NET941 NET949 NET905 NET947 NET928 NET951 
+ NET889 NET858 RE_RD1 RE_RD2 SAEB_RD1 SAEB_RD2 VDDHD VDDI VSSI WE_RD1 WE_RD2 
+ YL_RD1[0] YL_RD1[1] YL_RD2[0] YL_RD2[1] Y_DN_RD1[0] Y_DN_RD1[1] Y_DN_RD1[2] 
+ Y_DN_RD1[3] Y_DN_RD1[4] Y_DN_RD1[5] Y_DN_RD1[6] Y_DN_RD1[7] Y_DN_RD2[0] 
+ Y_DN_RD2[1] Y_DN_RD2[2] Y_DN_RD2[3] Y_DN_RD2[4] Y_DN_RD2[5] Y_DN_RD2[6] 
+ Y_DN_RD2[7] Y_UP_RD1[0] Y_UP_RD1[1] Y_UP_RD1[2] Y_UP_RD1[3] Y_UP_RD1[4] 
+ Y_UP_RD1[5] Y_UP_RD1[6] Y_UP_RD1[7] Y_UP_RD2[0] Y_UP_RD2[1] Y_UP_RD2[2] 
+ Y_UP_RD2[3] Y_UP_RD2[4] Y_UP_RD2[5] Y_UP_RD2[6] Y_UP_RD2[7] S1AHSF400W40_ARR_LIO_SIM
XARR_LIO_LDL BLB_LL_3 BLB_DUM_LL_3 NET0444[0] NET0444[1] NET0444[2] NET0444[3] 
+ NET0444[4] NET0444[5] NET0444[6] NET0444[7] NET0444[8] NET0444[9] 
+ NET0444[10] NET0444[11] NET0444[12] NET0444[13] BLB_LL_4 BLB_DUM_LL_4 
+ NET0446[0] NET0446[1] NET0446[2] NET0446[3] NET0446[4] NET0446[5] NET0446[6] 
+ NET0446[7] NET0446[8] NET0446[9] NET0446[10] NET0446[11] NET0446[12] 
+ NET0446[13] BLEQ_DN_LD4 BLEQ_DN_LD3 BLEQ_UP_LD4 BLEQ_UP_LD3 BL_LL_3 
+ BL_DUM_LL_3 NET0449[0] NET0449[1] NET0449[2] NET0449[3] NET0449[4] 
+ NET0449[5] NET0449[6] NET0449[7] NET0449[8] NET0449[9] NET0449[10] 
+ NET0449[11] NET0449[12] NET0449[13] BL_LL_4 BL_DUM_LL_4 NET0447[0] 
+ NET0447[1] NET0447[2] NET0447[3] NET0447[4] NET0447[5] NET0447[6] NET0447[7] 
+ NET0447[8] NET0447[9] NET0447[10] NET0447[11] NET0447[12] NET0447[13] VDDI 
+ GBLB_LL_3 GBLB_LL_4 GBL_LL_3 GBL_LL_4 GWB_LL_3 GWB_LL_4 GW_LL_3 GW_LL_4 
+ RE_LD4 RE_LD3 SAEB_LD4 SAEB_LD3 VDDHD VDDI VSSI WE_LD4 WE_LD3 YL_LD4[0] 
+ YL_LD4[1] YL_LD3[0] YL_LD3[1] Y_DN_LD4[0] Y_DN_LD4[1] Y_DN_LD4[2] 
+ Y_DN_LD4[3] Y_DN_LD4[4] Y_DN_LD4[5] Y_DN_LD4[6] Y_DN_LD4[7] Y_DN_LD3[0] 
+ Y_DN_LD3[1] Y_DN_LD3[2] Y_DN_LD3[3] Y_DN_LD3[4] Y_DN_LD3[5] Y_DN_LD3[6] 
+ Y_DN_LD3[7] Y_UP_LD4[0] Y_UP_LD4[1] Y_UP_LD4[2] Y_UP_LD4[3] Y_UP_LD4[4] 
+ Y_UP_LD4[5] Y_UP_LD4[6] Y_UP_LD4[7] Y_UP_LD3[0] Y_UP_LD3[1] Y_UP_LD3[2] 
+ Y_UP_LD3[3] Y_UP_LD3[4] Y_UP_LD3[5] Y_UP_LD3[6] Y_UP_LD3[7] S1AHSF400W40_ARR_LIO_SIM
XARR_MCB_RUR NET0928 NET0931 NET0929 NET0930 VDDI NET0926 NET0927 NET0925 
+ NET0918 VDDHD VDDI VSSI WL_RU3[0] WL_RU3[1] WL_RU4[0] WL_RU4[1] S1AHSF400W40_ARR_MCB_SIM
XARR_MCB_RUL NET0532 NET0910 NET0908 NET0911 VDDI NET0915 NET0914 NET0912 
+ NET0907 VDDHD VDDI VSSI WL_RU1[0] WL_RU1[1] WL_RU2[0] WL_RU2[1] S1AHSF400W40_ARR_MCB_SIM
XARR_MCB_LUR BL_LR_7 BL_DUM_LR_7 BLB_LR_7 BLB_DUM_LR_7 VDDI GBL_LR_78 
+ GBLB_LR_78 GW_LR_78 GWB_LR_78 VDDHD VDDI VSSI WL_LU2[0] WL_LU2[1] WL_LU1[0] 
+ WL_LU1[1] S1AHSF400W40_ARR_MCB_SIM
XARR_MCB_LDL BL_LL_2 BL_DUM_LL_2 BLB_LL_2 BLB_DUM_LL_2 VDDI GBL_LL_12 
+ GBLB_LL_12 GW_LL_12 GWB_LL_12 VDDHD VDDI VSSI WL_LD4[0] WL_LD4[1] WL_LD3[0] 
+ WL_LD3[1] S1AHSF400W40_ARR_MCB_SIM
XARR_MCB_RDR NET0941 NET0942 NET0940 NET0943 VDDI NET0947 NET0946 NET0944 
+ NET0945 VDDHD VDDI VSSI WL_RD3[0] WL_RD3[1] WL_RD4[0] WL_RD4[1] S1AHSF400W40_ARR_MCB_SIM
XARR_MCB_LDR BL_LR_2 BL_DUM_LR_2 BLB_LR_2 BLB_DUM_LR_2 VDDI GBL_LR_12 
+ GBLB_LR_12 GW_LR_12 GWB_LR_12 VDDHD VDDI VSSI WL_LD2[0] WL_LD2[1] WL_LD1[0] 
+ WL_LD1[1] S1AHSF400W40_ARR_MCB_SIM
XARR_MCB_LUL BL_LL_7 BL_DUM_LL_7 BLB_LL_7 BLB_DUM_LL_7 VDDI GBL_LL_78 
+ GBLB_LL_78 GW_LL_78 GWB_LL_78 VDDHD VDDI VSSI WL_LU4[0] WL_LU4[1] WL_LU3[0] 
+ WL_LU3[1] S1AHSF400W40_ARR_MCB_SIM
XARR_MCB_RDL NET0958 NET0957 NET0959 NET0956 VDDI NET0960 NET0961 NET0963 
+ NET0962 VDDHD VDDI VSSI WL_RD1[0] WL_RD1[1] WL_RD2[0] WL_RD2[1] S1AHSF400W40_ARR_MCB_SIM
XARR_WLLD_LU VDDI VDDHD VDDI VSSI WL_LU3[0] WL_LU3[1] WL_LU2[0] WL_LU2[1] 
+ S1AHSF400W40_ARR_WLLD_SIM
XARR_WLLD_RU VDDI VDDHD VDDI VSSI WL_RU2[0] WL_RU2[1] WL_RU3[0] WL_RU3[1] 
+ S1AHSF400W40_ARR_WLLD_SIM
XARR_WLLD_LD VDDI VDDHD VDDI VSSI WL_LD3[0] WL_LD3[1] WL_LD2[0] WL_LD2[1] 
+ S1AHSF400W40_ARR_WLLD_SIM
XARR_WLLD_RD VDDI VDDHD VDDI VSSI WL_RD2[0] WL_RD2[1] WL_RD3[0] WL_RD3[1] 
+ S1AHSF400W40_ARR_WLLD_SIM
XARR_BLLD_LUL BLB_LL_4 BLB_DUM_LL_4 BLB_LL_7 BLB_DUM_LL_7 BL_LL_4 BL_DUM_LL_4 
+ BL_LL_7 BL_DUM_LL_7 VDDI GBLB_LL_4 GBLB_LL_78 GBL_LL_4 GBL_LL_78 GWB_LL_4 
+ GWB_LL_78 GW_LL_4 GW_LL_78 VDDHD VDDI VSSI S1AHSF400W40_ARR_BLLD_SIM
XARRLBLLD_LDL BLB_LL_2 BLB_DUM_LL_2 BLB_LL_3 BLB_DUM_LL_3 BL_LL_2 BL_DUM_LL_2 
+ BL_LL_3 BL_DUM_LL_3 VDDI GBLB_LL_12 GBLB_LL_3 GBL_LL_12 GBL_LL_3 GWB_LL_12 
+ GWB_LL_3 GW_LL_12 GW_LL_3 VDDHD VDDI VSSI S1AHSF400W40_ARR_BLLD_SIM
XARR_BLLD_LDR BLB_LR_2 BLB_DUM_LR_2 BLB_LR_3 BLB_DUM_LR_3 BL_LR_2 BL_DUM_LR_2 
+ BL_LR_3 BL_DUM_LR_3 VDDI GBLB_LR_12 GBLB_LR_3 GBL_LR_12 GBL_LR_3 GWB_LR_12 
+ GWB_LR_3 GW_LR_12 GW_LR_3 VDDHD VDDI VSSI S1AHSF400W40_ARR_BLLD_SIM
XARR_BLLD_LUR BLB_LR_4 BLB_DUM_LR_4 BLB_LR_7 BLB_DUM_LR_7 BL_LR_4 BL_DUM_LR_4 
+ BL_LR_7 BL_DUM_LR_7 VDDI GBLB_LR_4 GBLB_LR_78 GBL_LR_4 GBL_LR_78 GWB_LR_4 
+ GWB_LR_78 GW_LR_4 GW_LR_78 VDDHD VDDI VSSI S1AHSF400W40_ARR_BLLD_SIM
XTKBL TRKBL BL_TK_TP VDDHD PD VDDHD VDDI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI WL_TK_ACT[0] 
+ WL_TK_ACT[1] WL_TK_ACT[2] WL_TK_ACT[3] WL_TK_ACT[4] WL_TK_ACT[5] 
+ WL_TK_ACT[6] WL_TK_ACT[7] WL_TK_ACT[8] WL_TK_ACT[9] WL_TK_ACT[10] 
+ WL_TK_ACT[11] WL_TK_ACT[12] WL_TK_ACT[13] WL_TK_ACT[14] WL_TK_ACT[15] 
+ WL_TK_ACT[16] WL_TK_ACT[17] WL_TK_ACT[18] WL_TK_ACT[19] WL_TK_ACT[20] 
+ WL_TK_ACT[21] WL_TK_ACT[22] WL_TK_ACT[23] WL_TK_ACT[24] WL_TK_ACT[25] 
+ WL_TK_ACT[26] WL_TK_ACT[27] WL_TK_ACT[28] WL_TK_ACT[29] WL_TK_ACT[30] 
+ WL_TK_ACT[31] WL_TK_ACT[32] WL_TK_ACT[33] WL_TK_ACT[34] WL_TK_ACT[35] 
+ WL_TK_ACT[36] WL_TK_ACT[37] WL_TK_ACT[38] WL_TK_ACT[39] WL_TK_ACT[40] 
+ WL_TK_ACT[41] WL_TK_ACT[42] WL_TK_ACT[43] WL_TK_ACT[44] WL_TK_ACT[45] 
+ WL_TK_ACT[46] WL_TK_ACT[47] WL_TK_ACT[48] WL_TK_ACT[49] WL_TK_ACT[50] 
+ WL_TK_ACT[51] WL_TK_ACT[52] WL_TK_ACT[53] WL_TK_ACT[54] WL_TK_ACT[55] 
+ WL_TK_ACT[56] WL_TK_ACT[57] WL_TK_ACT[58] WL_TK_ACT[59] WL_TK_ACT[60] 
+ WL_TK_ACT[61] WL_TK_ACT[62] WL_TK_ACT[63] WL_TK_ACT[64] WL_TK_ACT[65] 
+ WL_TK_ACT[66] WL_TK_ACT[67] WL_TK_ACT[68] WL_TK_ACT[69] WL_TK_ACT[70] 
+ WL_TK_ACT[71] WL_TK_ACT[72] WL_TK_ACT[73] WL_TK_ACT[74] WL_TK_ACT[75] 
+ WL_TK_ACT[76] WL_TK_ACT[77] WL_TK_ACT[78] WL_TK_ACT[79] WL_TK_ACT[80] 
+ WL_TK_ACT[81] WL_TK_ACT[82] WL_TK_ACT[83] WL_TK_ACT[84] WL_TK_ACT[85] 
+ WL_TK_ACT[86] WL_TK_ACT[87] WL_TK_ACT[88] WL_TK_ACT[89] WL_TK_ACT[90] 
+ WL_TK_ACT[91] WL_TK_ACT[92] WL_TK_ACT[93] WL_TK_ACT[94] WL_TK_ACT[95] 
+ WL_TK_ACT[96] WL_TK_ACT[97] WL_TK_ACT[98] WL_TK_ACT[99] WL_TK_ACT[100] 
+ WL_TK_ACT[101] WL_TK_ACT[102] WL_TK_ACT[103] WL_TK_ACT[104] WL_TK_ACT[105] 
+ WL_TK_ACT[106] WL_TK_ACT[107] WL_TK_ACT[108] WL_TK_ACT[109] WL_TK_ACT[110] 
+ WL_TK_ACT[111] WL_TK_ACT[112] WL_TK_ACT[113] WL_TK_ACT[114] WL_TK_ACT[115] 
+ WL_TK_ACT[116] WL_TK_ACT[117] WL_TK_ACT[118] WL_TK_ACT[119] WL_TK_ACT[120] 
+ WL_TK_ACT[121] WL_TK_ACT[122] WL_TK_ACT[123] WL_TK_ACT[124] WL_TK_ACT[125] 
+ WL_TK_ACT[126] WL_TK_ACT[127] WL_TK_ACT[128] WL_TK_ACT[129] WL_TK_ACT[130] 
+ WL_TK_ACT[131] WL_TK_ACT[132] WL_TK_ACT[133] WL_TK_ACT[134] WL_TK_ACT[135] 
+ WL_TK_ACT[136] WL_TK_ACT[137] WL_TK_ACT[138] WL_TK_ACT[139] WL_TK_ACT[140] 
+ WL_TK_ACT[141] WL_TK_ACT[142] WL_TK_ACT[143] WL_TK_ACT[144] WL_TK_ACT[145] 
+ WL_TK_ACT[146] WL_TK_ACT[147] WL_TK_ACT[148] WL_TK_ACT[149] WL_TK_ACT[150] 
+ WL_TK_ACT[151] WL_TK_ACT[152] WL_TK_ACT[153] WL_TK_ACT[154] WL_TK_ACT[155] 
+ WL_TK_ACT[156] WL_TK_ACT[157] WL_TK_ACT[158] WL_TK_ACT[159] WL_TK_ACT[160] 
+ WL_TK_ACT[161] WL_TK_ACT[162] WL_TK_ACT[163] WL_TK_ACT[164] WL_TK_ACT[165] 
+ WL_TK_ACT[166] WL_TK_ACT[167] WL_TK_ACT[168] WL_TK_ACT[169] WL_TK_ACT[170] 
+ WL_TK_ACT[171] WL_TK_ACT[172] WL_TK_ACT[173] WL_TK_ACT[174] WL_TK_ACT[175] 
+ WL_TK_ACT[176] WL_TK_ACT[177] WL_TK_ACT[178] WL_TK_ACT[179] WL_TK_ACT[180] 
+ WL_TK_ACT[181] WL_TK_ACT[182] WL_TK_ACT[183] WL_TK_ACT[184] WL_TK_ACT[185] 
+ WL_TK_ACT[186] WL_TK_ACT[187] WL_TK_ACT[188] WL_TK_ACT[189] WL_TK_ACT[190] 
+ WL_TK_ACT[191] WL_TK_ACT[192] WL_TK_ACT[193] WL_TK_ACT[194] WL_TK_ACT[195] 
+ WL_TK_ACT[196] WL_TK_ACT[197] WL_TK_ACT[198] WL_TK_ACT[199] WL_TK_ACT[200] 
+ WL_TK_ACT[201] WL_TK_ACT[202] WL_TK_ACT[203] WL_TK_ACT[204] WL_TK_ACT[205] 
+ WL_TK_ACT[206] WL_TK_ACT[207] WL_TK_ACT[208] WL_TK_ACT[209] WL_TK_ACT[210] 
+ WL_TK_ACT[211] WL_TK_ACT[212] WL_TK_ACT[213] WL_TK_ACT[214] WL_TK_ACT[215] 
+ WL_TK_ACT[216] WL_TK_ACT[217] WL_TK_ACT[218] WL_TK_ACT[219] WL_TK_ACT[220] 
+ WL_TK_ACT[221] WL_TK_ACT[222] WL_TK_ACT[223] WL_TK_ACT[224] WL_TK_ACT[225] 
+ WL_TK_ACT[226] WL_TK_ACT[227] WL_TK_ACT[228] WL_TK_ACT[229] WL_TK_ACT[230] 
+ WL_TK_ACT[231] WL_TK_ACT[232] WL_TK_ACT[233] WL_TK_ACT[234] WL_TK_ACT[235] 
+ WL_TK_ACT[236] WL_TK_ACT[237] WL_TK_ACT[238] WL_TK_ACT[239] WL_TK_ACT[240] 
+ WL_TK_ACT[241] WL_TK_ACT[242] WL_TK_ACT[243] WL_TK_ACT[244] WL_TK_ACT[245] 
+ WL_TK_ACT[246] WL_TK_ACT[247] WL_TK_ACT[248] WL_TK_ACT[249] WL_TK_ACT[250] 
+ WL_TK_ACT[251] WL_TK_ACT[252] WL_TK_ACT[253] WL_TK_ACT[254] WL_TK_ACT[255] 
+ WL_TK_ACT[256] WL_TK_ACT[257] WL_TK_ACT[258] WL_TK_ACT[259] WL_TK_ACT[260] 
+ WL_TK_ACT[261] WL_TK_ACT[262] WL_TK_ACT[263] WL_TK_ACT[264] WL_TK_ACT[265] 
+ WL_TK_ACT[266] WL_TK_ACT[267] WL_TK_ACT[268] WL_TK_ACT[269] WL_TK_ACT[270] 
+ WL_TK_ACT[271] WL_TK_ACT[272] WL_TK_ACT[273] WL_TK_ACT[274] WL_TK_ACT[275] 
+ WL_TK_ACT[276] WL_TK_ACT[277] WL_TK_ACT[278] WL_TK_ACT[279] WL_TK_ACT[280] 
+ WL_TK_ACT[281] WL_TK_ACT[282] WL_TK_ACT[283] WL_TK_ACT[284] WL_TK_ACT[285] 
+ WL_TK_ACT[286] WL_TK_ACT[287] WL_TK_ACT[288] WL_TK_ACT[289] WL_TK_ACT[290] 
+ WL_TK_ACT[291] WL_TK_ACT[292] WL_TK_ACT[293] WL_TK_ACT[294] WL_TK_ACT[295] 
+ WL_TK_ACT[296] WL_TK_ACT[297] WL_TK_ACT[298] WL_TK_ACT[299] WL_TK_ACT[300] 
+ WL_TK_ACT[301] WL_TK_ACT[302] WL_TK_ACT[303] WL_TK_ACT[304] WL_TK_ACT[305] 
+ WL_TK_ACT[306] WL_TK_ACT[307] WL_TK_ACT[308] WL_TK_ACT[309] WL_TK_ACT[310] 
+ WL_TK_ACT[311] WL_TK_ACT[312] WL_TK_ACT[313] WL_TK_ACT[314] WL_TK_ACT[315] 
+ WL_TK_ACT[316] WL_TK_ACT[317] WL_TK_ACT[318] WL_TK_ACT[319] WL_TK_ACT[320] 
+ WL_TK_ACT[321] WL_TK_ACT[322] WL_TK_ACT[323] WL_TK_ACT[324] WL_TK_ACT[325] 
+ WL_TK_ACT[326] WL_TK_ACT[327] WL_TK_ACT[328] WL_TK_ACT[329] WL_TK_ACT[330] 
+ WL_TK_ACT[331] WL_TK_ACT[332] WL_TK_ACT[333] WL_TK_ACT[334] WL_TK_ACT[335] 
+ WL_TK_ACT[336] WL_TK_ACT[337] WL_TK_ACT[338] WL_TK_ACT[339] WL_TK_ACT[340] 
+ WL_TK_ACT[341] WL_TK_ACT[342] WL_TK_ACT[343] WL_TK_ACT[344] WL_TK_ACT[345] 
+ WL_TK_ACT[346] WL_TK_ACT[347] WL_TK_ACT[348] WL_TK_ACT[349] WL_TK_ACT[350] 
+ WL_TK_ACT[351] WL_TK_ACT[352] WL_TK_ACT[353] WL_TK_ACT[354] WL_TK_ACT[355] 
+ WL_TK_ACT[356] WL_TK_ACT[357] WL_TK_ACT[358] WL_TK_ACT[359] WL_TK_ACT[360] 
+ WL_TK_ACT[361] WL_TK_ACT[362] WL_TK_ACT[363] WL_TK_ACT[364] WL_TK_ACT[365] 
+ WL_TK_ACT[366] WL_TK_ACT[367] WL_TK_ACT[368] WL_TK_ACT[369] WL_TK_ACT[370] 
+ WL_TK_ACT[371] WL_TK_ACT[372] WL_TK_ACT[373] WL_TK_ACT[374] WL_TK_ACT[375] 
+ WL_TK_ACT[376] WL_TK_ACT[377] WL_TK_ACT[378] WL_TK_ACT[379] WL_TK_ACT[380] 
+ WL_TK_ACT[381] WL_TK_ACT[382] WL_TK_ACT[383] WL_TK_ACT[384] WL_TK_ACT[385] 
+ WL_TK_ACT[386] WL_TK_ACT[387] WL_TK_ACT[388] WL_TK_ACT[389] WL_TK_ACT[390] 
+ WL_TK_ACT[391] WL_TK_ACT[392] WL_TK_ACT[393] WL_TK_ACT[394] WL_TK_ACT[395] 
+ WL_TK_ACT[396] WL_TK_ACT[397] WL_TK_ACT[398] WL_TK_ACT[399] WL_TK_ACT[400] 
+ WL_TK_ACT[401] WL_TK_ACT[402] WL_TK_ACT[403] WL_TK_ACT[404] WL_TK_ACT[405] 
+ WL_TK_ACT[406] WL_TK_ACT[407] WL_TK_ACT[408] WL_TK_ACT[409] WL_TK_ACT[410] 
+ WL_TK_ACT[411] WL_TK_ACT[412] WL_TK_ACT[413] WL_TK_ACT[414] WL_TK_ACT[415] 
+ WL_TK_ACT[416] WL_TK_ACT[417] WL_TK_ACT[418] WL_TK_ACT[419] WL_TK_ACT[420] 
+ WL_TK_ACT[421] WL_TK_ACT[422] WL_TK_ACT[423] WL_TK_ACT[424] WL_TK_ACT[425] 
+ WL_TK_ACT[426] WL_TK_ACT[427] WL_TK_ACT[428] WL_TK_ACT[429] WL_TK_ACT[430] 
+ WL_TK_ACT[431] WL_TK_ACT[432] WL_TK_ACT[433] WL_TK_ACT[434] WL_TK_ACT[435] 
+ WL_TK_ACT[436] WL_TK_ACT[437] WL_TK_ACT[438] WL_TK_ACT[439] WL_TK_ACT[440] 
+ WL_TK_ACT[441] WL_TK_ACT[442] WL_TK_ACT[443] WL_TK_ACT[444] WL_TK_ACT[445] 
+ WL_TK_ACT[446] WL_TK_ACT[447] WL_TK_ACT[448] WL_TK_ACT[449] WL_TK_ACT[450] 
+ WL_TK_ACT[451] WL_TK_ACT[452] WL_TK_ACT[453] WL_TK_ACT[454] WL_TK_ACT[455] 
+ WL_TK_ACT[456] WL_TK_ACT[457] WL_TK_ACT[458] WL_TK_ACT[459] WL_TK_ACT[460] 
+ WL_TK_ACT[461] WL_TK_ACT[462] WL_TK_ACT[463] WL_TK_ACT[464] WL_TK_ACT[465] 
+ WL_TK_ACT[466] WL_TK_ACT[467] WL_TK_ACT[468] WL_TK_ACT[469] WL_TK_ACT[470] 
+ WL_TK_ACT[471] WL_TK_ACT[472] WL_TK_ACT[473] WL_TK_ACT[474] WL_TK_ACT[475] 
+ WL_TK_ACT[476] WL_TK_ACT[477] WL_TK_ACT[478] WL_TK_ACT[479] WL_TK_ACT[480] 
+ WL_TK_ACT[481] WL_TK_ACT[482] WL_TK_ACT[483] WL_TK_ACT[484] WL_TK_ACT[485] 
+ WL_TK_ACT[486] WL_TK_ACT[487] WL_TK_ACT[488] WL_TK_ACT[489] WL_TK_ACT[490] 
+ WL_TK_ACT[491] WL_TK_ACT[492] WL_TK_ACT[493] WL_TK_ACT[494] WL_TK_ACT[495] 
+ WL_TK_ACT[496] WL_TK_ACT[497] WL_TK_ACT[498] WL_TK_ACT[499] WL_TK_ACT[500] 
+ WL_TK_ACT[501] WL_TK_ACT[502] WL_TK_ACT[503] WL_TK_ACT[504] WL_TK_ACT[505] 
+ WL_TK_ACT[506] WL_TK_ACT[507] WL_TK_ACT[508] WL_TK_ACT[509] WL_TK_ACT[510] 
+ WL_TK_ACT[511] TIEH_BT TIEL S1AHSF400W40_TKBL_SIM
XTKWL_LD VDDI TK_R2 TK_R3 VSSI WL_DUM_R2 WL_DUM_R3 WL_TK_R2 WL_TK_R3 
+ S1AHSF400W40_TKWL_LD_SIM
XTKWL_L VDDI TK TK_R2 VSSI WL_DUM_LT WL_DUM_R2 WL_TK WL_TK_R2 S1AHSF400W40_TKWL_SIM
XTKWL_R VDDI TK_R3 NET826 VSSI WL_DUM_R3 NET652 WL_TK_R3 WL_TK_LD S1AHSF400W40_TKWL_SIM
XIO_RL AWT2_L1 AWT2_R2 BIST2IO_L1 BIST2IO_R2 NET834 NET833 CKD_L1 CKD_R2 
+ NET836 NET837 NET827 NET830 NET832 NET831 PD_BUF_1 PD_BUF_R2 NET838 VDDHD 
+ VDDI VSSI WLP_SAEB_L1 WLP_SAEB_R2 S1AHSF400W40_IO_SIM
XIO_LR AWT2_L2 AWT2_L1 BIST2IO_L2 BIST2IO_L1 BWEBM_LR BWEB_LR CKD_L2 CKD_L1 
+ DM_LR D_LR GBLB_LR_12 GBL_LR_12 GWB_LR_12 GW_LR_12 PD_BUF_L2 PD_BUF_1 Q_LR 
+ VDDHD VDDI VSSI WLP_SAEB_L2 WLP_SAEB_L1 S1AHSF400W40_IO_SIM
XIO_LL AWT2_L4 AWT2_L3 BIST2IO_L4 BIST2IO_L3 BWEBM_LL BWEB_LL CKD_L4 CKD_L3 
+ DM_LL D_LL GBLB_LL_12 GBL_LL_12 GWB_LL_12 GW_LL_12 PD_BUF_L4 PD_BUF_L3 Q_LL 
+ VDDHD VDDI VSSI WLP_SAEB_L4 WLP_SAEB_L3 S1AHSF400W40_IO_SIM
XIO_RR AWT2_R3 AWT2_R4 BIST2IO_R3 BIST2IO_R4 NET847 NET848 CKD_R3 CKD_R4 
+ NET846 NET844 NET855 NET854 NET850 NET853 PD_BUF_R3 PD_BUF_R4 NET843 VDDHD 
+ VDDI VSSI WLP_SAEB_R3 WLP_SAEB_R4 S1AHSF400W40_IO_SIM
XIO_LD_L AWT2_L3 AWT2_L2 BIST2IO_L3 BIST2IO_L2 CKD_L3 CKD_L2 PD_BUF_L3 
+ PD_BUF_L2 VDDHD VDDI VSSI WLP_SAEB_L3 WLP_SAEB_L2 S1AHSF400W40_IO_LD_SIM
XIO_LD_R AWT2_R2 AWT2_R3 BIST2IO_R2 BIST2IO_R3 CKD_R2 CKD_R3 PD_BUF_R2 
+ PD_BUF_R3 VDDHD VDDI VSSI WLP_SAEB_R2 WLP_SAEB_R3 S1AHSF400W40_IO_LD_SIM
XCNT AWT AWT2_L1 BIST BIST2IO_L1 WL_TK CEB CEBM CKD_L1 CLK VDDHD VDDI 
+ DEC_X0_1[0] DEC_X0_1[1] DEC_X0_1[2] DEC_X0_1[3] DEC_X0_1[4] DEC_X0_1[5] 
+ DEC_X0_1[6] DEC_X0_1[7] DEC_X1_1[0] DEC_X1_1[1] DEC_X1_1[2] DEC_X1_1[3] 
+ DEC_X1_1[4] DEC_X1_1[5] DEC_X1_1[6] DEC_X1_1[7] DEC_X2_1[0] DEC_X2_1[1] 
+ DEC_X2_1[2] DEC_X2_1[3] DEC_X3_1[0] DEC_X3_1[1] DEC_X3_1[2] DEC_X3_1[3] 
+ DEC_X3_1[4] DEC_X3_1[5] DEC_X3_1[6] DEC_X3_1[7] DEC_Y_1[0] DEC_Y_1[1] 
+ DEC_Y_1[2] DEC_Y_1[3] DEC_Y_1[4] DEC_Y_1[5] DEC_Y_1[6] DEC_Y_1[7] FAD1[0] 
+ FAD1[1] FAD1[2] FAD1[3] FAD1[4] FAD1[5] FAD1[6] FAD1[7] FAD1[8] FAD1[9] 
+ FAD1[10] FAD2[0] FAD2[1] FAD2[2] FAD2[3] FAD2[4] FAD2[5] FAD2[6] FAD2[7] 
+ FAD2[8] FAD2[9] FAD2[10] NET934[0] NET934[1] PD PD_BUF_1 PD_CVDDBUF_1 PTSEL 
+ REDEN_BT REDEN1 REDEN2 REDENB_BT RSTB RTSEL[0] RTSEL[1] RW_RE_1 SCLK SDIN 
+ SDOUT TK TM TRKBL VDDHD VDDI VHI_LT VLO_LT VSSI WEB WEBM WLP_SAE_1 
+ WLP_SAEB_L1 WLP_SAE_TK_1 WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] 
+ X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] 
+ XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL_1[0] YM[0] YM[1] YM[2] YM[3] 
+ S1AHSF400W40_CNT_SIM
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_STRAP_888_U_386
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_STRAP_888_U_386 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_X2_SHARE PD_BUF VDDHD 
+ VDDI VSSI
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2[4]:B DEC_X2[5]:B DEC_X2[6]:B DEC_X2[7]:B DEC_X2_SHARE:B 
*.PININFO PD_BUF:B VDDHD:B VDDI:B VSSI:B
XSTRAP DEC_X2[6] DEC_X2_SHARE VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_888_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_STRAP_888_U_384
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_STRAP_888_U_384 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_X2_SHARE PD_BUF VDDHD 
+ VDDI VSSI
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2[4]:B DEC_X2[5]:B DEC_X2[6]:B DEC_X2[7]:B DEC_X2_SHARE:B 
*.PININFO PD_BUF:B VDDHD:B VDDI:B VSSI:B
XSTRAP DEC_X2[5] DEC_X2_SHARE VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_888_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_STRAP_882_U_66
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_STRAP_882_U_66 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2_SHARE 
+ PD_BUF VDDHD VDDI VSSI
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2_SHARE:B PD_BUF:B VDDHD:B 
*.PININFO VDDI:B VSSI:B
XSTRAP DEC_X2[1] DEC_X2_SHARE VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_882_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_STRAP_882_U_128
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_STRAP_882_U_128 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2_SHARE 
+ PD_BUF VDDHD VDDI VSSI
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2_SHARE:B PD_BUF:B VDDHD:B 
*.PININFO VDDI:B VSSI:B
XSTRAP DEC_X2[1] DEC_X2_SHARE VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_882_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_STRAP_888_U_258
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_STRAP_888_U_258 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_X2_SHARE PD_BUF VDDHD 
+ VDDI VSSI
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2[4]:B DEC_X2[5]:B DEC_X2[6]:B DEC_X2[7]:B DEC_X2_SHARE:B 
*.PININFO PD_BUF:B VDDHD:B VDDI:B VSSI:B
XSTRAP DEC_X2[4] DEC_X2_SHARE VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_888_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_STRAP_884_U_130
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_STRAP_884_U_130 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2_SHARE:B PD_BUF:B VDDHD:B VDDI:B VSSI:B
XSTRAP DEC_X2[2] DEC_X2_SHARE VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_884_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_STRAP_884_U_256
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_STRAP_884_U_256 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2_SHARE PD_BUF VDDHD VDDI VSSI
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2_SHARE:B PD_BUF:B VDDHD:B VDDI:B VSSI:B
XSTRAP DEC_X2[3] DEC_X2_SHARE VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_884_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_STRAP_888_U_512
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_STRAP_888_U_512 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_X2_SHARE PD_BUF VDDHD 
+ VDDI VSSI
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2[4]:B DEC_X2[5]:B DEC_X2[6]:B DEC_X2[7]:B DEC_X2_SHARE:B 
*.PININFO PD_BUF:B VDDHD:B VDDI:B VSSI:B
XSTRAP DEC_X2[7] DEC_X2_SHARE VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_888_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_STRAP_U_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_STRAP_U_SIM DEC_X0_BT[0] DEC_X0_BT[1] DEC_X0_BT[2] DEC_X0_BT[3] 
+ DEC_X0_BT[4] DEC_X0_BT[5] DEC_X0_BT[6] DEC_X0_BT[7] DEC_X0_TP[0] 
+ DEC_X0_TP[1] DEC_X0_TP[2] DEC_X0_TP[3] DEC_X0_TP[4] DEC_X0_TP[5] 
+ DEC_X0_TP[6] DEC_X0_TP[7] DEC_X1_BT[0] DEC_X1_BT[1] DEC_X1_BT[2] 
+ DEC_X1_BT[3] DEC_X1_BT[4] DEC_X1_BT[5] DEC_X1_BT[6] DEC_X1_BT[7] 
+ DEC_X1_TP[0] DEC_X1_TP[1] DEC_X1_TP[2] DEC_X1_TP[3] DEC_X1_TP[4] 
+ DEC_X1_TP[5] DEC_X1_TP[6] DEC_X1_TP[7] DEC_X2_BT[0] DEC_X2_BT[1] 
+ DEC_X2_BT[2] DEC_X2_BT[3] DEC_X2_BT[4] DEC_X2_BT[5] DEC_X2_BT[6] 
+ DEC_X2_BT[7] DEC_X2_SHARE DEC_X2_TP[0] DEC_X2_TP[1] DEC_X2_TP[2] 
+ DEC_X2_TP[3] DEC_X2_TP[4] DEC_X2_TP[5] DEC_X2_TP[6] DEC_X2_TP[7] PD_BUF_BT 
+ PD_BUF_TP VDDHD VDDI VSSI
*.PININFO DEC_X0_BT[0]:I DEC_X0_BT[1]:I DEC_X0_BT[2]:I DEC_X0_BT[3]:I 
*.PININFO DEC_X0_BT[4]:I DEC_X0_BT[5]:I DEC_X0_BT[6]:I DEC_X0_BT[7]:I 
*.PININFO DEC_X1_BT[0]:I DEC_X1_BT[1]:I DEC_X1_BT[2]:I DEC_X1_BT[3]:I 
*.PININFO DEC_X1_BT[4]:I DEC_X1_BT[5]:I DEC_X1_BT[6]:I DEC_X1_BT[7]:I 
*.PININFO PD_BUF_BT:I DEC_X0_TP[0]:O DEC_X0_TP[1]:O DEC_X0_TP[2]:O 
*.PININFO DEC_X0_TP[3]:O DEC_X0_TP[4]:O DEC_X0_TP[5]:O DEC_X0_TP[6]:O 
*.PININFO DEC_X0_TP[7]:O DEC_X1_TP[0]:O DEC_X1_TP[1]:O DEC_X1_TP[2]:O 
*.PININFO DEC_X1_TP[3]:O DEC_X1_TP[4]:O DEC_X1_TP[5]:O DEC_X1_TP[6]:O 
*.PININFO DEC_X1_TP[7]:O PD_BUF_TP:O DEC_X2_BT[0]:B DEC_X2_BT[1]:B 
*.PININFO DEC_X2_BT[2]:B DEC_X2_BT[3]:B DEC_X2_BT[4]:B DEC_X2_BT[5]:B 
*.PININFO DEC_X2_BT[6]:B DEC_X2_BT[7]:B DEC_X2_SHARE:B DEC_X2_TP[0]:B 
*.PININFO DEC_X2_TP[1]:B DEC_X2_TP[2]:B DEC_X2_TP[3]:B DEC_X2_TP[4]:B 
*.PININFO DEC_X2_TP[5]:B DEC_X2_TP[6]:B DEC_X2_TP[7]:B VDDHD:B VDDI:B VSSI:B
XI32 NET064[0] NET064[1] NET064[2] NET064[3] NET064[4] NET064[5] NET064[6] 
+ NET064[7] NET062[0] NET062[1] NET062[2] NET062[3] NET062[4] NET062[5] 
+ NET062[6] NET062[7] NET063[0] NET063[1] NET063[2] NET063[3] NET063[4] 
+ NET063[5] NET063[6] NET063[7] NET065 NET058 NET061 NET060 NET059 
+ S1AHSF400W40_SB_STRAP_888_U_386
XI33 NET072[0] NET072[1] NET072[2] NET072[3] NET072[4] NET072[5] NET072[6] 
+ NET072[7] NET070[0] NET070[1] NET070[2] NET070[3] NET070[4] NET070[5] 
+ NET070[6] NET070[7] NET071[0] NET071[1] NET071[2] NET071[3] NET071[4] 
+ NET071[5] NET071[6] NET071[7] NET073 NET066 NET069 NET068 NET067 
+ S1AHSF400W40_SB_STRAP_888_U_384
XI31 NET079[0] NET079[1] NET079[2] NET079[3] NET079[4] NET079[5] NET079[6] 
+ NET079[7] NET080[0] NET080[1] NET080[2] NET080[3] NET080[4] NET080[5] 
+ NET080[6] NET080[7] NET078[0] NET078[1] NET081 NET074 NET077 NET076 NET075 
+ S1AHSF400W40_SB_STRAP_882_U_66
XI26 NET025[0] NET025[1] NET025[2] NET025[3] NET025[4] NET025[5] NET025[6] 
+ NET025[7] NET044[0] NET044[1] NET044[2] NET044[3] NET044[4] NET044[5] 
+ NET044[6] NET044[7] NET046[0] NET046[1] NET026 NET01 NET08 NET02 NET06 
+ S1AHSF400W40_SB_STRAP_882_U_128
XI30 NET014[0] NET014[1] NET014[2] NET014[3] NET014[4] NET014[5] NET014[6] 
+ NET014[7] NET07[0] NET07[1] NET07[2] NET07[3] NET07[4] NET07[5] NET07[6] 
+ NET07[7] NET015[0] NET015[1] NET015[2] NET015[3] NET015[4] NET015[5] 
+ NET015[6] NET015[7] NET013 NET017 NET024 NET040 NET011 S1AHSF400W40_SB_STRAP_888_U_258
XI29 NET041[0] NET041[1] NET041[2] NET041[3] NET041[4] NET041[5] NET041[6] 
+ NET041[7] NET039[0] NET039[1] NET039[2] NET039[3] NET039[4] NET039[5] 
+ NET039[6] NET039[7] NET038[0] NET038[1] NET038[2] NET038[3] NET018 NET037 
+ NET012 NET010 NET016 S1AHSF400W40_SB_STRAP_884_U_130
XI27 NET027[0] NET027[1] NET027[2] NET027[3] NET027[4] NET027[5] NET027[6] 
+ NET027[7] NET03[0] NET03[1] NET03[2] NET03[3] NET03[4] NET03[5] NET03[6] 
+ NET03[7] NET09[0] NET09[1] NET09[2] NET09[3] NET028 NET021 NET05 NET023 
+ NET022 S1AHSF400W40_SB_STRAP_884_U_256
XI28 NET035[0] NET035[1] NET035[2] NET035[3] NET035[4] NET035[5] NET035[6] 
+ NET035[7] NET033[0] NET033[1] NET033[2] NET033[3] NET033[4] NET033[5] 
+ NET033[6] NET033[7] NET034[0] NET034[1] NET034[2] NET034[3] NET034[4] 
+ NET034[5] NET034[6] NET034[7] NET036 NET029 NET032 NET031 NET030 
+ S1AHSF400W40_SB_STRAP_888_U_512
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_888_LD_D_384
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_888_LD_D_384 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_X2_SHARE[0] PD_BUF 
+ VDDHD VDDI VSSI
*.PININFO PD_BUF:I DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2[4]:B DEC_X2[5]:B DEC_X2[6]:B DEC_X2[7]:B DEC_X2_SHARE[0]:B 
*.PININFO VDDHD:B VDDI:B VSSI:B
XI171<1> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2_SHARE[0] PD_BUF VDDHD VDDI VSSI 
+ NET027[0] NET027[1] NET027[2] NET027[3] NET027[4] NET027[5] NET027[6] 
+ NET027[7] NET027[8] NET027[9] NET027[10] NET027[11] NET027[12] NET027[13] 
+ NET027[14] NET027[15] NET027[16] NET027[17] NET027[18] NET027[19] NET027[20] 
+ NET027[21] NET027[22] NET027[23] NET027[24] NET027[25] NET027[26] NET027[27] 
+ NET027[28] NET027[29] NET027[30] NET027[31] NET027[32] NET027[33] NET027[34] 
+ NET027[35] NET027[36] NET027[37] NET027[38] NET027[39] NET027[40] NET027[41] 
+ NET027[42] NET027[43] NET027[44] NET027[45] NET027[46] NET027[47] NET027[48] 
+ NET027[49] NET027[50] NET027[51] NET027[52] NET027[53] NET027[54] NET027[55] 
+ NET027[56] NET027[57] NET027[58] NET027[59] NET027[60] NET027[61] NET027[62] 
+ NET027[63] S1AHSF400W40_WLDV_64X1_888_SB
XWLDV<4> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[4] DEC_X2_SHARE[4] PD_BUF VDDHD VDDI VSSI 
+ NET40[0] NET40[1] NET40[2] NET40[3] NET40[4] NET40[5] NET40[6] NET40[7] 
+ NET40[8] NET40[9] NET40[10] NET40[11] NET40[12] NET40[13] NET40[14] 
+ NET40[15] NET40[16] NET40[17] NET40[18] NET40[19] NET40[20] NET40[21] 
+ NET40[22] NET40[23] NET40[24] NET40[25] NET40[26] NET40[27] NET40[28] 
+ NET40[29] NET40[30] NET40[31] NET40[32] NET40[33] NET40[34] NET40[35] 
+ NET40[36] NET40[37] NET40[38] NET40[39] NET40[40] NET40[41] NET40[42] 
+ NET40[43] NET40[44] NET40[45] NET40[46] NET40[47] NET40[48] NET40[49] 
+ NET40[50] NET40[51] NET40[52] NET40[53] NET40[54] NET40[55] NET40[56] 
+ NET40[57] NET40[58] NET40[59] NET40[60] NET40[61] NET40[62] NET40[63] 
+ S1AHSF400W40_WLDV_64X1_888_SB
XWLDV_64X1<3> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[3] DEC_X2_SHARE[3] PD_BUF VDDHD VDDI 
+ VSSI NET58[0] NET58[1] NET58[2] NET58[3] NET58[4] NET58[5] NET58[6] NET58[7] 
+ NET58[8] NET58[9] NET58[10] NET58[11] NET58[12] NET58[13] NET58[14] 
+ NET58[15] NET58[16] NET58[17] NET58[18] NET58[19] NET58[20] NET58[21] 
+ NET58[22] NET58[23] NET58[24] NET58[25] NET58[26] NET58[27] NET58[28] 
+ NET58[29] NET58[30] NET58[31] NET58[32] NET58[33] NET58[34] NET58[35] 
+ NET58[36] NET58[37] NET58[38] NET58[39] NET58[40] NET58[41] NET58[42] 
+ NET58[43] NET58[44] NET58[45] NET58[46] NET58[47] NET58[48] NET58[49] 
+ NET58[50] NET58[51] NET58[52] NET58[53] NET58[54] NET58[55] NET58[56] 
+ NET58[57] NET58[58] NET58[59] NET58[60] NET58[61] NET58[62] NET58[63] 
+ S1AHSF400W40_WLDV_64X1_888_SB
XWLDV_64X1<1> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[1] DEC_X2_SHARE[1] PD_BUF VDDHD VDDI 
+ VSSI NET67[0] NET67[1] NET67[2] NET67[3] NET67[4] NET67[5] NET67[6] NET67[7] 
+ NET67[8] NET67[9] NET67[10] NET67[11] NET67[12] NET67[13] NET67[14] 
+ NET67[15] NET67[16] NET67[17] NET67[18] NET67[19] NET67[20] NET67[21] 
+ NET67[22] NET67[23] NET67[24] NET67[25] NET67[26] NET67[27] NET67[28] 
+ NET67[29] NET67[30] NET67[31] NET67[32] NET67[33] NET67[34] NET67[35] 
+ NET67[36] NET67[37] NET67[38] NET67[39] NET67[40] NET67[41] NET67[42] 
+ NET67[43] NET67[44] NET67[45] NET67[46] NET67[47] NET67[48] NET67[49] 
+ NET67[50] NET67[51] NET67[52] NET67[53] NET67[54] NET67[55] NET67[56] 
+ NET67[57] NET67[58] NET67[59] NET67[60] NET67[61] NET67[62] NET67[63] 
+ S1AHSF400W40_WLDV_64X1_888_SB
XWLDV_64X1<2> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[2] DEC_X2_SHARE[2] PD_BUF VDDHD VDDI 
+ VSSI NET76[0] NET76[1] NET76[2] NET76[3] NET76[4] NET76[5] NET76[6] NET76[7] 
+ NET76[8] NET76[9] NET76[10] NET76[11] NET76[12] NET76[13] NET76[14] 
+ NET76[15] NET76[16] NET76[17] NET76[18] NET76[19] NET76[20] NET76[21] 
+ NET76[22] NET76[23] NET76[24] NET76[25] NET76[26] NET76[27] NET76[28] 
+ NET76[29] NET76[30] NET76[31] NET76[32] NET76[33] NET76[34] NET76[35] 
+ NET76[36] NET76[37] NET76[38] NET76[39] NET76[40] NET76[41] NET76[42] 
+ NET76[43] NET76[44] NET76[45] NET76[46] NET76[47] NET76[48] NET76[49] 
+ NET76[50] NET76[51] NET76[52] NET76[53] NET76[54] NET76[55] NET76[56] 
+ NET76[57] NET76[58] NET76[59] NET76[60] NET76[61] NET76[62] NET76[63] 
+ S1AHSF400W40_WLDV_64X1_888_SB
XI160 DEC_X2[4] DEC_X2_SHARE[4] VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_888_SB
XSTRAP2 DEC_X2[2] DEC_X2_SHARE[2] VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_888_SB
XSTRAP1 DEC_X2[1] DEC_X2_SHARE[1] VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_888_SB
XSTRAP3 DEC_X2[3] DEC_X2_SHARE[3] VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_888_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_888_LD_D_386
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_888_LD_D_386 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_X2_SHARE[0] PD_BUF 
+ VDDHD VDDI VSSI
*.PININFO PD_BUF:I DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2[4]:B DEC_X2[5]:B DEC_X2[6]:B DEC_X2[7]:B DEC_X2_SHARE[0]:B 
*.PININFO VDDHD:B VDDI:B VSSI:B
XI171<1> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2_SHARE[0] PD_BUF VDDHD VDDI VSSI 
+ NET027[0] NET027[1] NET027[2] NET027[3] NET027[4] NET027[5] NET027[6] 
+ NET027[7] NET027[8] NET027[9] NET027[10] NET027[11] NET027[12] NET027[13] 
+ NET027[14] NET027[15] NET027[16] NET027[17] NET027[18] NET027[19] NET027[20] 
+ NET027[21] NET027[22] NET027[23] NET027[24] NET027[25] NET027[26] NET027[27] 
+ NET027[28] NET027[29] NET027[30] NET027[31] NET027[32] NET027[33] NET027[34] 
+ NET027[35] NET027[36] NET027[37] NET027[38] NET027[39] NET027[40] NET027[41] 
+ NET027[42] NET027[43] NET027[44] NET027[45] NET027[46] NET027[47] NET027[48] 
+ NET027[49] NET027[50] NET027[51] NET027[52] NET027[53] NET027[54] NET027[55] 
+ NET027[56] NET027[57] NET027[58] NET027[59] NET027[60] NET027[61] NET027[62] 
+ NET027[63] S1AHSF400W40_WLDV_64X1_888_SB
XWLDV<4> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[4] DEC_X2_SHARE[4] PD_BUF VDDHD VDDI VSSI 
+ NET40[0] NET40[1] NET40[2] NET40[3] NET40[4] NET40[5] NET40[6] NET40[7] 
+ NET40[8] NET40[9] NET40[10] NET40[11] NET40[12] NET40[13] NET40[14] 
+ NET40[15] NET40[16] NET40[17] NET40[18] NET40[19] NET40[20] NET40[21] 
+ NET40[22] NET40[23] NET40[24] NET40[25] NET40[26] NET40[27] NET40[28] 
+ NET40[29] NET40[30] NET40[31] NET40[32] NET40[33] NET40[34] NET40[35] 
+ NET40[36] NET40[37] NET40[38] NET40[39] NET40[40] NET40[41] NET40[42] 
+ NET40[43] NET40[44] NET40[45] NET40[46] NET40[47] NET40[48] NET40[49] 
+ NET40[50] NET40[51] NET40[52] NET40[53] NET40[54] NET40[55] NET40[56] 
+ NET40[57] NET40[58] NET40[59] NET40[60] NET40[61] NET40[62] NET40[63] 
+ S1AHSF400W40_WLDV_64X1_888_SB
XWLDV_64X1<3> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[3] DEC_X2_SHARE[3] PD_BUF VDDHD VDDI 
+ VSSI NET58[0] NET58[1] NET58[2] NET58[3] NET58[4] NET58[5] NET58[6] NET58[7] 
+ NET58[8] NET58[9] NET58[10] NET58[11] NET58[12] NET58[13] NET58[14] 
+ NET58[15] NET58[16] NET58[17] NET58[18] NET58[19] NET58[20] NET58[21] 
+ NET58[22] NET58[23] NET58[24] NET58[25] NET58[26] NET58[27] NET58[28] 
+ NET58[29] NET58[30] NET58[31] NET58[32] NET58[33] NET58[34] NET58[35] 
+ NET58[36] NET58[37] NET58[38] NET58[39] NET58[40] NET58[41] NET58[42] 
+ NET58[43] NET58[44] NET58[45] NET58[46] NET58[47] NET58[48] NET58[49] 
+ NET58[50] NET58[51] NET58[52] NET58[53] NET58[54] NET58[55] NET58[56] 
+ NET58[57] NET58[58] NET58[59] NET58[60] NET58[61] NET58[62] NET58[63] 
+ S1AHSF400W40_WLDV_64X1_888_SB
XWLDV_64X1<1> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[1] DEC_X2_SHARE[1] PD_BUF VDDHD VDDI 
+ VSSI NET67[0] NET67[1] NET67[2] NET67[3] NET67[4] NET67[5] NET67[6] NET67[7] 
+ NET67[8] NET67[9] NET67[10] NET67[11] NET67[12] NET67[13] NET67[14] 
+ NET67[15] NET67[16] NET67[17] NET67[18] NET67[19] NET67[20] NET67[21] 
+ NET67[22] NET67[23] NET67[24] NET67[25] NET67[26] NET67[27] NET67[28] 
+ NET67[29] NET67[30] NET67[31] NET67[32] NET67[33] NET67[34] NET67[35] 
+ NET67[36] NET67[37] NET67[38] NET67[39] NET67[40] NET67[41] NET67[42] 
+ NET67[43] NET67[44] NET67[45] NET67[46] NET67[47] NET67[48] NET67[49] 
+ NET67[50] NET67[51] NET67[52] NET67[53] NET67[54] NET67[55] NET67[56] 
+ NET67[57] NET67[58] NET67[59] NET67[60] NET67[61] NET67[62] NET67[63] 
+ S1AHSF400W40_WLDV_64X1_888_SB
XWLDV_64X1<2> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[2] DEC_X2_SHARE[2] PD_BUF VDDHD VDDI 
+ VSSI NET76[0] NET76[1] NET76[2] NET76[3] NET76[4] NET76[5] NET76[6] NET76[7] 
+ NET76[8] NET76[9] NET76[10] NET76[11] NET76[12] NET76[13] NET76[14] 
+ NET76[15] NET76[16] NET76[17] NET76[18] NET76[19] NET76[20] NET76[21] 
+ NET76[22] NET76[23] NET76[24] NET76[25] NET76[26] NET76[27] NET76[28] 
+ NET76[29] NET76[30] NET76[31] NET76[32] NET76[33] NET76[34] NET76[35] 
+ NET76[36] NET76[37] NET76[38] NET76[39] NET76[40] NET76[41] NET76[42] 
+ NET76[43] NET76[44] NET76[45] NET76[46] NET76[47] NET76[48] NET76[49] 
+ NET76[50] NET76[51] NET76[52] NET76[53] NET76[54] NET76[55] NET76[56] 
+ NET76[57] NET76[58] NET76[59] NET76[60] NET76[61] NET76[62] NET76[63] 
+ S1AHSF400W40_WLDV_64X1_888_SB
XI160 DEC_X2[4] DEC_X2_SHARE[4] VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_888_SB
XSTRAP2 DEC_X2[2] DEC_X2_SHARE[2] VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_888_SB
XSTRAP1 DEC_X2[1] DEC_X2_SHARE[1] VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_888_SB
XSTRAP3 DEC_X2[3] DEC_X2_SHARE[3] VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_888_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_882_LD_D_66
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_882_LD_D_66 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2_SHARE[0] 
+ PD_BUF VDDHD VDDI VSSI
*.PININFO PD_BUF:I DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2_SHARE[0]:B VDDHD:B VDDI:B 
*.PININFO VSSI:B
XWLDV_64X1<0> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2_SHARE[0] PD_BUF VDDHD VDDI 
+ VSSI NET18[0] NET18[1] NET18[2] NET18[3] NET18[4] NET18[5] NET18[6] NET18[7] 
+ NET18[8] NET18[9] NET18[10] NET18[11] NET18[12] NET18[13] NET18[14] 
+ NET18[15] NET18[16] NET18[17] NET18[18] NET18[19] NET18[20] NET18[21] 
+ NET18[22] NET18[23] NET18[24] NET18[25] NET18[26] NET18[27] NET18[28] 
+ NET18[29] NET18[30] NET18[31] NET18[32] NET18[33] NET18[34] NET18[35] 
+ NET18[36] NET18[37] NET18[38] NET18[39] NET18[40] NET18[41] NET18[42] 
+ NET18[43] NET18[44] NET18[45] NET18[46] NET18[47] NET18[48] NET18[49] 
+ NET18[50] NET18[51] NET18[52] NET18[53] NET18[54] NET18[55] NET18[56] 
+ NET18[57] NET18[58] NET18[59] NET18[60] NET18[61] NET18[62] NET18[63] 
+ S1AHSF400W40_WLDV_64X1_882_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_882_LD_D_128
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_882_LD_D_128 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2_SHARE[0] 
+ PD_BUF VDDHD VDDI VSSI
*.PININFO PD_BUF:I DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2_SHARE[0]:B VDDHD:B VDDI:B 
*.PININFO VSSI:B
XI171<1> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2_SHARE[0] PD_BUF VDDHD VDDI VSSI 
+ NET18[0] NET18[1] NET18[2] NET18[3] NET18[4] NET18[5] NET18[6] NET18[7] 
+ NET18[8] NET18[9] NET18[10] NET18[11] NET18[12] NET18[13] NET18[14] 
+ NET18[15] NET18[16] NET18[17] NET18[18] NET18[19] NET18[20] NET18[21] 
+ NET18[22] NET18[23] NET18[24] NET18[25] NET18[26] NET18[27] NET18[28] 
+ NET18[29] NET18[30] NET18[31] NET18[32] NET18[33] NET18[34] NET18[35] 
+ NET18[36] NET18[37] NET18[38] NET18[39] NET18[40] NET18[41] NET18[42] 
+ NET18[43] NET18[44] NET18[45] NET18[46] NET18[47] NET18[48] NET18[49] 
+ NET18[50] NET18[51] NET18[52] NET18[53] NET18[54] NET18[55] NET18[56] 
+ NET18[57] NET18[58] NET18[59] NET18[60] NET18[61] NET18[62] NET18[63] 
+ S1AHSF400W40_WLDV_64X1_882_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_884_LD_D_130
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_884_LD_D_130 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2_SHARE[0] PD_BUF VDDHD VDDI VSSI
*.PININFO PD_BUF:I DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2_SHARE[0]:B VDDHD:B VDDI:B VSSI:B
XWLDV_64X1<0> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2_SHARE[0] PD_BUF VDDHD VDDI 
+ VSSI NET027[0] NET027[1] NET027[2] NET027[3] NET027[4] NET027[5] NET027[6] 
+ NET027[7] NET027[8] NET027[9] NET027[10] NET027[11] NET027[12] NET027[13] 
+ NET027[14] NET027[15] NET027[16] NET027[17] NET027[18] NET027[19] NET027[20] 
+ NET027[21] NET027[22] NET027[23] NET027[24] NET027[25] NET027[26] NET027[27] 
+ NET027[28] NET027[29] NET027[30] NET027[31] NET027[32] NET027[33] NET027[34] 
+ NET027[35] NET027[36] NET027[37] NET027[38] NET027[39] NET027[40] NET027[41] 
+ NET027[42] NET027[43] NET027[44] NET027[45] NET027[46] NET027[47] NET027[48] 
+ NET027[49] NET027[50] NET027[51] NET027[52] NET027[53] NET027[54] NET027[55] 
+ NET027[56] NET027[57] NET027[58] NET027[59] NET027[60] NET027[61] NET027[62] 
+ NET027[63] S1AHSF400W40_WLDV_64X1_884_SB
XWLDV_64X1<1> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[1] DEC_X2_SHARE[1] PD_BUF VDDHD VDDI 
+ VSSI NET67[0] NET67[1] NET67[2] NET67[3] NET67[4] NET67[5] NET67[6] NET67[7] 
+ NET67[8] NET67[9] NET67[10] NET67[11] NET67[12] NET67[13] NET67[14] 
+ NET67[15] NET67[16] NET67[17] NET67[18] NET67[19] NET67[20] NET67[21] 
+ NET67[22] NET67[23] NET67[24] NET67[25] NET67[26] NET67[27] NET67[28] 
+ NET67[29] NET67[30] NET67[31] NET67[32] NET67[33] NET67[34] NET67[35] 
+ NET67[36] NET67[37] NET67[38] NET67[39] NET67[40] NET67[41] NET67[42] 
+ NET67[43] NET67[44] NET67[45] NET67[46] NET67[47] NET67[48] NET67[49] 
+ NET67[50] NET67[51] NET67[52] NET67[53] NET67[54] NET67[55] NET67[56] 
+ NET67[57] NET67[58] NET67[59] NET67[60] NET67[61] NET67[62] NET67[63] 
+ S1AHSF400W40_WLDV_64X1_884_SB
XSTRAP1 DEC_X2[1] DEC_X2_SHARE[1] VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_884_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_888_LD_D_258
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_888_LD_D_258 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_X2_SHARE[0] PD_BUF 
+ VDDHD VDDI VSSI
*.PININFO PD_BUF:I DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2[4]:B DEC_X2[5]:B DEC_X2[6]:B DEC_X2[7]:B DEC_X2_SHARE[0]:B 
*.PININFO VDDHD:B VDDI:B VSSI:B
XI171<1> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2_SHARE[0] PD_BUF VDDHD VDDI VSSI 
+ NET027[0] NET027[1] NET027[2] NET027[3] NET027[4] NET027[5] NET027[6] 
+ NET027[7] NET027[8] NET027[9] NET027[10] NET027[11] NET027[12] NET027[13] 
+ NET027[14] NET027[15] NET027[16] NET027[17] NET027[18] NET027[19] NET027[20] 
+ NET027[21] NET027[22] NET027[23] NET027[24] NET027[25] NET027[26] NET027[27] 
+ NET027[28] NET027[29] NET027[30] NET027[31] NET027[32] NET027[33] NET027[34] 
+ NET027[35] NET027[36] NET027[37] NET027[38] NET027[39] NET027[40] NET027[41] 
+ NET027[42] NET027[43] NET027[44] NET027[45] NET027[46] NET027[47] NET027[48] 
+ NET027[49] NET027[50] NET027[51] NET027[52] NET027[53] NET027[54] NET027[55] 
+ NET027[56] NET027[57] NET027[58] NET027[59] NET027[60] NET027[61] NET027[62] 
+ NET027[63] S1AHSF400W40_WLDV_64X1_888_SB
XWLDV_64X1<1> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[1] DEC_X2_SHARE[1] PD_BUF VDDHD VDDI 
+ VSSI NET67[0] NET67[1] NET67[2] NET67[3] NET67[4] NET67[5] NET67[6] NET67[7] 
+ NET67[8] NET67[9] NET67[10] NET67[11] NET67[12] NET67[13] NET67[14] 
+ NET67[15] NET67[16] NET67[17] NET67[18] NET67[19] NET67[20] NET67[21] 
+ NET67[22] NET67[23] NET67[24] NET67[25] NET67[26] NET67[27] NET67[28] 
+ NET67[29] NET67[30] NET67[31] NET67[32] NET67[33] NET67[34] NET67[35] 
+ NET67[36] NET67[37] NET67[38] NET67[39] NET67[40] NET67[41] NET67[42] 
+ NET67[43] NET67[44] NET67[45] NET67[46] NET67[47] NET67[48] NET67[49] 
+ NET67[50] NET67[51] NET67[52] NET67[53] NET67[54] NET67[55] NET67[56] 
+ NET67[57] NET67[58] NET67[59] NET67[60] NET67[61] NET67[62] NET67[63] 
+ S1AHSF400W40_WLDV_64X1_888_SB
XWLDV_64X1<2> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[2] DEC_X2_SHARE[2] PD_BUF VDDHD VDDI 
+ VSSI NET76[0] NET76[1] NET76[2] NET76[3] NET76[4] NET76[5] NET76[6] NET76[7] 
+ NET76[8] NET76[9] NET76[10] NET76[11] NET76[12] NET76[13] NET76[14] 
+ NET76[15] NET76[16] NET76[17] NET76[18] NET76[19] NET76[20] NET76[21] 
+ NET76[22] NET76[23] NET76[24] NET76[25] NET76[26] NET76[27] NET76[28] 
+ NET76[29] NET76[30] NET76[31] NET76[32] NET76[33] NET76[34] NET76[35] 
+ NET76[36] NET76[37] NET76[38] NET76[39] NET76[40] NET76[41] NET76[42] 
+ NET76[43] NET76[44] NET76[45] NET76[46] NET76[47] NET76[48] NET76[49] 
+ NET76[50] NET76[51] NET76[52] NET76[53] NET76[54] NET76[55] NET76[56] 
+ NET76[57] NET76[58] NET76[59] NET76[60] NET76[61] NET76[62] NET76[63] 
+ S1AHSF400W40_WLDV_64X1_888_SB
XSTRAP2 DEC_X2[2] DEC_X2_SHARE[2] VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_888_SB
XSTRAP1 DEC_X2[1] DEC_X2_SHARE[1] VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_888_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_884_LD_D_256
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_884_LD_D_256 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2_SHARE[0] PD_BUF VDDHD VDDI VSSI
*.PININFO PD_BUF:I DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2_SHARE[0]:B VDDHD:B VDDI:B VSSI:B
XWLDV_64X1<0> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2_SHARE[0] PD_BUF VDDHD VDDI 
+ VSSI NET027[0] NET027[1] NET027[2] NET027[3] NET027[4] NET027[5] NET027[6] 
+ NET027[7] NET027[8] NET027[9] NET027[10] NET027[11] NET027[12] NET027[13] 
+ NET027[14] NET027[15] NET027[16] NET027[17] NET027[18] NET027[19] NET027[20] 
+ NET027[21] NET027[22] NET027[23] NET027[24] NET027[25] NET027[26] NET027[27] 
+ NET027[28] NET027[29] NET027[30] NET027[31] NET027[32] NET027[33] NET027[34] 
+ NET027[35] NET027[36] NET027[37] NET027[38] NET027[39] NET027[40] NET027[41] 
+ NET027[42] NET027[43] NET027[44] NET027[45] NET027[46] NET027[47] NET027[48] 
+ NET027[49] NET027[50] NET027[51] NET027[52] NET027[53] NET027[54] NET027[55] 
+ NET027[56] NET027[57] NET027[58] NET027[59] NET027[60] NET027[61] NET027[62] 
+ NET027[63] S1AHSF400W40_WLDV_64X1_884_SB
XWLDV_64X1<1> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[1] DEC_X2_SHARE[1] PD_BUF VDDHD VDDI 
+ VSSI NET67[0] NET67[1] NET67[2] NET67[3] NET67[4] NET67[5] NET67[6] NET67[7] 
+ NET67[8] NET67[9] NET67[10] NET67[11] NET67[12] NET67[13] NET67[14] 
+ NET67[15] NET67[16] NET67[17] NET67[18] NET67[19] NET67[20] NET67[21] 
+ NET67[22] NET67[23] NET67[24] NET67[25] NET67[26] NET67[27] NET67[28] 
+ NET67[29] NET67[30] NET67[31] NET67[32] NET67[33] NET67[34] NET67[35] 
+ NET67[36] NET67[37] NET67[38] NET67[39] NET67[40] NET67[41] NET67[42] 
+ NET67[43] NET67[44] NET67[45] NET67[46] NET67[47] NET67[48] NET67[49] 
+ NET67[50] NET67[51] NET67[52] NET67[53] NET67[54] NET67[55] NET67[56] 
+ NET67[57] NET67[58] NET67[59] NET67[60] NET67[61] NET67[62] NET67[63] 
+ S1AHSF400W40_WLDV_64X1_884_SB
XWLDV_64X1<2> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[2] DEC_X2_SHARE[2] PD_BUF VDDHD VDDI 
+ VSSI NET76[0] NET76[1] NET76[2] NET76[3] NET76[4] NET76[5] NET76[6] NET76[7] 
+ NET76[8] NET76[9] NET76[10] NET76[11] NET76[12] NET76[13] NET76[14] 
+ NET76[15] NET76[16] NET76[17] NET76[18] NET76[19] NET76[20] NET76[21] 
+ NET76[22] NET76[23] NET76[24] NET76[25] NET76[26] NET76[27] NET76[28] 
+ NET76[29] NET76[30] NET76[31] NET76[32] NET76[33] NET76[34] NET76[35] 
+ NET76[36] NET76[37] NET76[38] NET76[39] NET76[40] NET76[41] NET76[42] 
+ NET76[43] NET76[44] NET76[45] NET76[46] NET76[47] NET76[48] NET76[49] 
+ NET76[50] NET76[51] NET76[52] NET76[53] NET76[54] NET76[55] NET76[56] 
+ NET76[57] NET76[58] NET76[59] NET76[60] NET76[61] NET76[62] NET76[63] 
+ S1AHSF400W40_WLDV_64X1_884_SB
XSTRAP2 DEC_X2[2] DEC_X2_SHARE[2] VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_884_SB
XSTRAP1 DEC_X2[1] DEC_X2_SHARE[1] VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_884_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_WLDV_888_LD_D_512
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_WLDV_888_LD_D_512 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] DEC_X2_SHARE[0] PD_BUF 
+ VDDHD VDDI VSSI
*.PININFO PD_BUF:I DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X2[4]:B DEC_X2[5]:B DEC_X2[6]:B DEC_X2[7]:B DEC_X2_SHARE[0]:B 
*.PININFO VDDHD:B VDDI:B VSSI:B
XI171<1> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2_SHARE[0] PD_BUF VDDHD VDDI VSSI 
+ NET027[0] NET027[1] NET027[2] NET027[3] NET027[4] NET027[5] NET027[6] 
+ NET027[7] NET027[8] NET027[9] NET027[10] NET027[11] NET027[12] NET027[13] 
+ NET027[14] NET027[15] NET027[16] NET027[17] NET027[18] NET027[19] NET027[20] 
+ NET027[21] NET027[22] NET027[23] NET027[24] NET027[25] NET027[26] NET027[27] 
+ NET027[28] NET027[29] NET027[30] NET027[31] NET027[32] NET027[33] NET027[34] 
+ NET027[35] NET027[36] NET027[37] NET027[38] NET027[39] NET027[40] NET027[41] 
+ NET027[42] NET027[43] NET027[44] NET027[45] NET027[46] NET027[47] NET027[48] 
+ NET027[49] NET027[50] NET027[51] NET027[52] NET027[53] NET027[54] NET027[55] 
+ NET027[56] NET027[57] NET027[58] NET027[59] NET027[60] NET027[61] NET027[62] 
+ NET027[63] S1AHSF400W40_WLDV_64X1_888_SB
XWLDV<4> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[4] DEC_X2_SHARE[4] PD_BUF VDDHD VDDI VSSI 
+ NET40[0] NET40[1] NET40[2] NET40[3] NET40[4] NET40[5] NET40[6] NET40[7] 
+ NET40[8] NET40[9] NET40[10] NET40[11] NET40[12] NET40[13] NET40[14] 
+ NET40[15] NET40[16] NET40[17] NET40[18] NET40[19] NET40[20] NET40[21] 
+ NET40[22] NET40[23] NET40[24] NET40[25] NET40[26] NET40[27] NET40[28] 
+ NET40[29] NET40[30] NET40[31] NET40[32] NET40[33] NET40[34] NET40[35] 
+ NET40[36] NET40[37] NET40[38] NET40[39] NET40[40] NET40[41] NET40[42] 
+ NET40[43] NET40[44] NET40[45] NET40[46] NET40[47] NET40[48] NET40[49] 
+ NET40[50] NET40[51] NET40[52] NET40[53] NET40[54] NET40[55] NET40[56] 
+ NET40[57] NET40[58] NET40[59] NET40[60] NET40[61] NET40[62] NET40[63] 
+ S1AHSF400W40_WLDV_64X1_888_SB
XWLDV_64X1<3> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[3] DEC_X2_SHARE[3] PD_BUF VDDHD VDDI 
+ VSSI NET58[0] NET58[1] NET58[2] NET58[3] NET58[4] NET58[5] NET58[6] NET58[7] 
+ NET58[8] NET58[9] NET58[10] NET58[11] NET58[12] NET58[13] NET58[14] 
+ NET58[15] NET58[16] NET58[17] NET58[18] NET58[19] NET58[20] NET58[21] 
+ NET58[22] NET58[23] NET58[24] NET58[25] NET58[26] NET58[27] NET58[28] 
+ NET58[29] NET58[30] NET58[31] NET58[32] NET58[33] NET58[34] NET58[35] 
+ NET58[36] NET58[37] NET58[38] NET58[39] NET58[40] NET58[41] NET58[42] 
+ NET58[43] NET58[44] NET58[45] NET58[46] NET58[47] NET58[48] NET58[49] 
+ NET58[50] NET58[51] NET58[52] NET58[53] NET58[54] NET58[55] NET58[56] 
+ NET58[57] NET58[58] NET58[59] NET58[60] NET58[61] NET58[62] NET58[63] 
+ S1AHSF400W40_WLDV_64X1_888_SB
XI158<3> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[5] DEC_X2_SHARE[5] PD_BUF VDDHD VDDI VSSI 
+ NET49[0] NET49[1] NET49[2] NET49[3] NET49[4] NET49[5] NET49[6] NET49[7] 
+ NET49[8] NET49[9] NET49[10] NET49[11] NET49[12] NET49[13] NET49[14] 
+ NET49[15] NET49[16] NET49[17] NET49[18] NET49[19] NET49[20] NET49[21] 
+ NET49[22] NET49[23] NET49[24] NET49[25] NET49[26] NET49[27] NET49[28] 
+ NET49[29] NET49[30] NET49[31] NET49[32] NET49[33] NET49[34] NET49[35] 
+ NET49[36] NET49[37] NET49[38] NET49[39] NET49[40] NET49[41] NET49[42] 
+ NET49[43] NET49[44] NET49[45] NET49[46] NET49[47] NET49[48] NET49[49] 
+ NET49[50] NET49[51] NET49[52] NET49[53] NET49[54] NET49[55] NET49[56] 
+ NET49[57] NET49[58] NET49[59] NET49[60] NET49[61] NET49[62] NET49[63] 
+ S1AHSF400W40_WLDV_64X1_888_SB
XWLDV_64X1<1> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[1] DEC_X2_SHARE[1] PD_BUF VDDHD VDDI 
+ VSSI NET67[0] NET67[1] NET67[2] NET67[3] NET67[4] NET67[5] NET67[6] NET67[7] 
+ NET67[8] NET67[9] NET67[10] NET67[11] NET67[12] NET67[13] NET67[14] 
+ NET67[15] NET67[16] NET67[17] NET67[18] NET67[19] NET67[20] NET67[21] 
+ NET67[22] NET67[23] NET67[24] NET67[25] NET67[26] NET67[27] NET67[28] 
+ NET67[29] NET67[30] NET67[31] NET67[32] NET67[33] NET67[34] NET67[35] 
+ NET67[36] NET67[37] NET67[38] NET67[39] NET67[40] NET67[41] NET67[42] 
+ NET67[43] NET67[44] NET67[45] NET67[46] NET67[47] NET67[48] NET67[49] 
+ NET67[50] NET67[51] NET67[52] NET67[53] NET67[54] NET67[55] NET67[56] 
+ NET67[57] NET67[58] NET67[59] NET67[60] NET67[61] NET67[62] NET67[63] 
+ S1AHSF400W40_WLDV_64X1_888_SB
XI163<3> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[6] DEC_X2_SHARE[6] PD_BUF VDDHD VDDI VSSI 
+ NET31[0] NET31[1] NET31[2] NET31[3] NET31[4] NET31[5] NET31[6] NET31[7] 
+ NET31[8] NET31[9] NET31[10] NET31[11] NET31[12] NET31[13] NET31[14] 
+ NET31[15] NET31[16] NET31[17] NET31[18] NET31[19] NET31[20] NET31[21] 
+ NET31[22] NET31[23] NET31[24] NET31[25] NET31[26] NET31[27] NET31[28] 
+ NET31[29] NET31[30] NET31[31] NET31[32] NET31[33] NET31[34] NET31[35] 
+ NET31[36] NET31[37] NET31[38] NET31[39] NET31[40] NET31[41] NET31[42] 
+ NET31[43] NET31[44] NET31[45] NET31[46] NET31[47] NET31[48] NET31[49] 
+ NET31[50] NET31[51] NET31[52] NET31[53] NET31[54] NET31[55] NET31[56] 
+ NET31[57] NET31[58] NET31[59] NET31[60] NET31[61] NET31[62] NET31[63] 
+ S1AHSF400W40_WLDV_64X1_888_SB
XWLDV_64X1<2> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[2] DEC_X2_SHARE[2] PD_BUF VDDHD VDDI 
+ VSSI NET76[0] NET76[1] NET76[2] NET76[3] NET76[4] NET76[5] NET76[6] NET76[7] 
+ NET76[8] NET76[9] NET76[10] NET76[11] NET76[12] NET76[13] NET76[14] 
+ NET76[15] NET76[16] NET76[17] NET76[18] NET76[19] NET76[20] NET76[21] 
+ NET76[22] NET76[23] NET76[24] NET76[25] NET76[26] NET76[27] NET76[28] 
+ NET76[29] NET76[30] NET76[31] NET76[32] NET76[33] NET76[34] NET76[35] 
+ NET76[36] NET76[37] NET76[38] NET76[39] NET76[40] NET76[41] NET76[42] 
+ NET76[43] NET76[44] NET76[45] NET76[46] NET76[47] NET76[48] NET76[49] 
+ NET76[50] NET76[51] NET76[52] NET76[53] NET76[54] NET76[55] NET76[56] 
+ NET76[57] NET76[58] NET76[59] NET76[60] NET76[61] NET76[62] NET76[63] 
+ S1AHSF400W40_WLDV_64X1_888_SB
XI160 DEC_X2[4] DEC_X2_SHARE[4] VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_888_SB
XI161 DEC_X2[5] DEC_X2_SHARE[5] VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_888_SB
XI162 DEC_X2[6] DEC_X2_SHARE[6] VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_888_SB
XSTRAP2 DEC_X2[2] DEC_X2_SHARE[2] VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_888_SB
XSTRAP1 DEC_X2[1] DEC_X2_SHARE[1] VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_888_SB
XSTRAP3 DEC_X2[3] DEC_X2_SHARE[3] VDDHD VDDI VSSI S1AHSF400W40_XDRV_STRAP_888_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SB_BK_LD_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SB_BK_LD_SIM DEC_X0_BT[0] DEC_X0_BT[1] DEC_X0_BT[2] DEC_X0_BT[3] 
+ DEC_X0_BT[4] DEC_X0_BT[5] DEC_X0_BT[6] DEC_X0_BT[7] DEC_X0_TP[0] 
+ DEC_X0_TP[1] DEC_X0_TP[2] DEC_X0_TP[3] DEC_X0_TP[4] DEC_X0_TP[5] 
+ DEC_X0_TP[6] DEC_X0_TP[7] DEC_X1_BT[0] DEC_X1_BT[1] DEC_X1_BT[2] 
+ DEC_X1_BT[3] DEC_X1_BT[4] DEC_X1_BT[5] DEC_X1_BT[6] DEC_X1_BT[7] 
+ DEC_X1_TP[0] DEC_X1_TP[1] DEC_X1_TP[2] DEC_X1_TP[3] DEC_X1_TP[4] 
+ DEC_X1_TP[5] DEC_X1_TP[6] DEC_X1_TP[7] DEC_X2_BT[0] DEC_X2_BT[1] 
+ DEC_X2_BT[2] DEC_X2_BT[3] DEC_X2_BT[4] DEC_X2_BT[5] DEC_X2_BT[6] 
+ DEC_X2_BT[7] DEC_X2_SHARE[0] DEC_X2_TP[0] DEC_X2_TP[1] DEC_X2_TP[2] 
+ DEC_X2_TP[3] DEC_X2_TP[4] DEC_X2_TP[5] DEC_X2_TP[6] DEC_X2_TP[7] PD_BUF_BT 
+ PD_BUF_TP VDDHD VDDI VSSI
*.PININFO DEC_X0_BT[0]:B DEC_X0_BT[1]:B DEC_X0_BT[2]:B DEC_X0_BT[3]:B 
*.PININFO DEC_X0_BT[4]:B DEC_X0_BT[5]:B DEC_X0_BT[6]:B DEC_X0_BT[7]:B 
*.PININFO DEC_X0_TP[0]:B DEC_X0_TP[1]:B DEC_X0_TP[2]:B DEC_X0_TP[3]:B 
*.PININFO DEC_X0_TP[4]:B DEC_X0_TP[5]:B DEC_X0_TP[6]:B DEC_X0_TP[7]:B 
*.PININFO DEC_X1_BT[0]:B DEC_X1_BT[1]:B DEC_X1_BT[2]:B DEC_X1_BT[3]:B 
*.PININFO DEC_X1_BT[4]:B DEC_X1_BT[5]:B DEC_X1_BT[6]:B DEC_X1_BT[7]:B 
*.PININFO DEC_X1_TP[0]:B DEC_X1_TP[1]:B DEC_X1_TP[2]:B DEC_X1_TP[3]:B 
*.PININFO DEC_X1_TP[4]:B DEC_X1_TP[5]:B DEC_X1_TP[6]:B DEC_X1_TP[7]:B 
*.PININFO DEC_X2_BT[0]:B DEC_X2_BT[1]:B DEC_X2_BT[2]:B DEC_X2_BT[3]:B 
*.PININFO DEC_X2_BT[4]:B DEC_X2_BT[5]:B DEC_X2_BT[6]:B DEC_X2_BT[7]:B 
*.PININFO DEC_X2_SHARE[0]:B DEC_X2_TP[0]:B DEC_X2_TP[1]:B DEC_X2_TP[2]:B 
*.PININFO DEC_X2_TP[3]:B DEC_X2_TP[4]:B DEC_X2_TP[5]:B DEC_X2_TP[6]:B 
*.PININFO DEC_X2_TP[7]:B PD_BUF_BT:B PD_BUF_TP:B VDDHD:B VDDI:B VSSI:B
XI34 NET012[0] NET012[1] NET012[2] NET012[3] NET012[4] NET012[5] NET012[6] 
+ NET012[7] NET049[0] NET049[1] NET049[2] NET049[3] NET049[4] NET049[5] 
+ NET049[6] NET049[7] NET061[0] NET061[1] NET061[2] NET061[3] NET061[4] 
+ NET061[5] NET061[6] NET061[7] NET043 NET062 NET057 NET053 NET019 
+ S1AHSF400W40_SB_WLDV_888_LD_D_384
XI33 NET048[0] NET048[1] NET048[2] NET048[3] NET048[4] NET048[5] NET048[6] 
+ NET048[7] NET064[0] NET064[1] NET064[2] NET064[3] NET064[4] NET064[5] 
+ NET064[6] NET064[7] NET063[0] NET063[1] NET063[2] NET063[3] NET063[4] 
+ NET063[5] NET063[6] NET063[7] NET046 NET058 NET04 NET045 NET042 
+ S1AHSF400W40_SB_WLDV_888_LD_D_386
XI32 NET039[0] NET039[1] NET039[2] NET039[3] NET039[4] NET039[5] NET039[6] 
+ NET039[7] NET037[0] NET037[1] NET037[2] NET037[3] NET037[4] NET037[5] 
+ NET037[6] NET037[7] NET060[0] NET060[1] NET038 NET052 NET056 NET065 NET066 
+ S1AHSF400W40_SB_WLDV_882_LD_D_66
XI28 NET020[0] NET020[1] NET020[2] NET020[3] NET020[4] NET020[5] NET020[6] 
+ NET020[7] NET018[0] NET018[1] NET018[2] NET018[3] NET018[4] NET018[5] 
+ NET018[6] NET018[7] NET017[0] NET017[1] NET059 NET01 NET016 NET014 NET015 
+ S1AHSF400W40_SB_WLDV_882_LD_D_128
XI30 NET06[0] NET06[1] NET06[2] NET06[3] NET06[4] NET06[5] NET06[6] NET06[7] 
+ NET011[0] NET011[1] NET011[2] NET011[3] NET011[4] NET011[5] NET011[6] 
+ NET011[7] NET010[0] NET010[1] NET010[2] NET010[3] NET09 NET07 NET03 NET02 
+ NET05 S1AHSF400W40_SB_WLDV_884_LD_D_130
XI29 NET08[0] NET08[1] NET08[2] NET08[3] NET08[4] NET08[5] NET08[6] NET08[7] 
+ NET028[0] NET028[1] NET028[2] NET028[3] NET028[4] NET028[5] NET028[6] 
+ NET028[7] NET023[0] NET023[1] NET023[2] NET023[3] NET023[4] NET023[5] 
+ NET023[6] NET023[7] NET027 NET022 NET026 NET024 NET025 S1AHSF400W40_SB_WLDV_888_LD_D_258
XI26 NET18[0] NET18[1] NET18[2] NET18[3] NET18[4] NET18[5] NET18[6] NET18[7] 
+ NET17[0] NET17[1] NET17[2] NET17[3] NET17[4] NET17[5] NET17[6] NET17[7] 
+ NET021[0] NET021[1] NET021[2] NET021[3] NET013 NET12 NET16 NET14 NET15 
+ S1AHSF400W40_SB_WLDV_884_LD_D_256
XI27 NET036[0] NET036[1] NET036[2] NET036[3] NET036[4] NET036[5] NET036[6] 
+ NET036[7] NET035[0] NET035[1] NET035[2] NET035[3] NET035[4] NET035[5] 
+ NET035[6] NET035[7] NET030[0] NET030[1] NET030[2] NET030[3] NET030[4] 
+ NET030[5] NET030[6] NET030[7] NET034 NET029 NET033 NET031 NET032 
+ S1AHSF400W40_SB_WLDV_888_LD_D_512
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SIM_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SIM_SB AWT BIST BWEBM_LL BWEBM_LR BWEB_LL BWEB_LR CEB CEBM CLK DM_LL 
+ DM_LR D_LL D_LR PD PTSEL Q_LL Q_LR RTSEL[0] RTSEL[1] TM VDDI VSSI WEB WEBM 
+ WL_TK_ACT[0] WL_TK_ACT[1] WL_TK_ACT[2] WL_TK_ACT[3] WL_TK_ACT[4] 
+ WL_TK_ACT[5] WL_TK_ACT[6] WL_TK_ACT[7] WL_TK_ACT[8] WL_TK_ACT[9] 
+ WL_TK_ACT[10] WL_TK_ACT[11] WL_TK_ACT[12] WL_TK_ACT[13] WL_TK_ACT[14] 
+ WL_TK_ACT[15] WL_TK_ACT[16] WL_TK_ACT[17] WL_TK_ACT[18] WL_TK_ACT[19] 
+ WL_TK_ACT[20] WL_TK_ACT[21] WL_TK_ACT[22] WL_TK_ACT[23] WL_TK_ACT[24] 
+ WL_TK_ACT[25] WL_TK_ACT[26] WL_TK_ACT[27] WL_TK_ACT[28] WL_TK_ACT[29] 
+ WL_TK_ACT[30] WL_TK_ACT[31] WL_TK_ACT[32] WL_TK_ACT[33] WL_TK_ACT[34] 
+ WL_TK_ACT[35] WL_TK_ACT[36] WL_TK_ACT[37] WL_TK_ACT[38] WL_TK_ACT[39] 
+ WL_TK_ACT[40] WL_TK_ACT[41] WL_TK_ACT[42] WL_TK_ACT[43] WL_TK_ACT[44] 
+ WL_TK_ACT[45] WL_TK_ACT[46] WL_TK_ACT[47] WL_TK_ACT[48] WL_TK_ACT[49] 
+ WL_TK_ACT[50] WL_TK_ACT[51] WL_TK_ACT[52] WL_TK_ACT[53] WL_TK_ACT[54] 
+ WL_TK_ACT[55] WL_TK_ACT[56] WL_TK_ACT[57] WL_TK_ACT[58] WL_TK_ACT[59] 
+ WL_TK_ACT[60] WL_TK_ACT[61] WL_TK_ACT[62] WL_TK_ACT[63] WL_TK_ACT[64] 
+ WL_TK_ACT[65] WL_TK_ACT[66] WL_TK_ACT[67] WL_TK_ACT[68] WL_TK_ACT[69] 
+ WL_TK_ACT[70] WL_TK_ACT[71] WL_TK_ACT[72] WL_TK_ACT[73] WL_TK_ACT[74] 
+ WL_TK_ACT[75] WL_TK_ACT[76] WL_TK_ACT[77] WL_TK_ACT[78] WL_TK_ACT[79] 
+ WL_TK_ACT[80] WL_TK_ACT[81] WL_TK_ACT[82] WL_TK_ACT[83] WL_TK_ACT[84] 
+ WL_TK_ACT[85] WL_TK_ACT[86] WL_TK_ACT[87] WL_TK_ACT[88] WL_TK_ACT[89] 
+ WL_TK_ACT[90] WL_TK_ACT[91] WL_TK_ACT[92] WL_TK_ACT[93] WL_TK_ACT[94] 
+ WL_TK_ACT[95] WL_TK_ACT[96] WL_TK_ACT[97] WL_TK_ACT[98] WL_TK_ACT[99] 
+ WL_TK_ACT[100] WL_TK_ACT[101] WL_TK_ACT[102] WL_TK_ACT[103] WL_TK_ACT[104] 
+ WL_TK_ACT[105] WL_TK_ACT[106] WL_TK_ACT[107] WL_TK_ACT[108] WL_TK_ACT[109] 
+ WL_TK_ACT[110] WL_TK_ACT[111] WL_TK_ACT[112] WL_TK_ACT[113] WL_TK_ACT[114] 
+ WL_TK_ACT[115] WL_TK_ACT[116] WL_TK_ACT[117] WL_TK_ACT[118] WL_TK_ACT[119] 
+ WL_TK_ACT[120] WL_TK_ACT[121] WL_TK_ACT[122] WL_TK_ACT[123] WL_TK_ACT[124] 
+ WL_TK_ACT[125] WL_TK_ACT[126] WL_TK_ACT[127] WL_TK_ACT[128] WL_TK_ACT[129] 
+ WL_TK_ACT[130] WL_TK_ACT[131] WL_TK_ACT[132] WL_TK_ACT[133] WL_TK_ACT[134] 
+ WL_TK_ACT[135] WL_TK_ACT[136] WL_TK_ACT[137] WL_TK_ACT[138] WL_TK_ACT[139] 
+ WL_TK_ACT[140] WL_TK_ACT[141] WL_TK_ACT[142] WL_TK_ACT[143] WL_TK_ACT[144] 
+ WL_TK_ACT[145] WL_TK_ACT[146] WL_TK_ACT[147] WL_TK_ACT[148] WL_TK_ACT[149] 
+ WL_TK_ACT[150] WL_TK_ACT[151] WL_TK_ACT[152] WL_TK_ACT[153] WL_TK_ACT[154] 
+ WL_TK_ACT[155] WL_TK_ACT[156] WL_TK_ACT[157] WL_TK_ACT[158] WL_TK_ACT[159] 
+ WL_TK_ACT[160] WL_TK_ACT[161] WL_TK_ACT[162] WL_TK_ACT[163] WL_TK_ACT[164] 
+ WL_TK_ACT[165] WL_TK_ACT[166] WL_TK_ACT[167] WL_TK_ACT[168] WL_TK_ACT[169] 
+ WL_TK_ACT[170] WL_TK_ACT[171] WL_TK_ACT[172] WL_TK_ACT[173] WL_TK_ACT[174] 
+ WL_TK_ACT[175] WL_TK_ACT[176] WL_TK_ACT[177] WL_TK_ACT[178] WL_TK_ACT[179] 
+ WL_TK_ACT[180] WL_TK_ACT[181] WL_TK_ACT[182] WL_TK_ACT[183] WL_TK_ACT[184] 
+ WL_TK_ACT[185] WL_TK_ACT[186] WL_TK_ACT[187] WL_TK_ACT[188] WL_TK_ACT[189] 
+ WL_TK_ACT[190] WL_TK_ACT[191] WL_TK_ACT[192] WL_TK_ACT[193] WL_TK_ACT[194] 
+ WL_TK_ACT[195] WL_TK_ACT[196] WL_TK_ACT[197] WL_TK_ACT[198] WL_TK_ACT[199] 
+ WL_TK_ACT[200] WL_TK_ACT[201] WL_TK_ACT[202] WL_TK_ACT[203] WL_TK_ACT[204] 
+ WL_TK_ACT[205] WL_TK_ACT[206] WL_TK_ACT[207] WL_TK_ACT[208] WL_TK_ACT[209] 
+ WL_TK_ACT[210] WL_TK_ACT[211] WL_TK_ACT[212] WL_TK_ACT[213] WL_TK_ACT[214] 
+ WL_TK_ACT[215] WL_TK_ACT[216] WL_TK_ACT[217] WL_TK_ACT[218] WL_TK_ACT[219] 
+ WL_TK_ACT[220] WL_TK_ACT[221] WL_TK_ACT[222] WL_TK_ACT[223] WL_TK_ACT[224] 
+ WL_TK_ACT[225] WL_TK_ACT[226] WL_TK_ACT[227] WL_TK_ACT[228] WL_TK_ACT[229] 
+ WL_TK_ACT[230] WL_TK_ACT[231] WL_TK_ACT[232] WL_TK_ACT[233] WL_TK_ACT[234] 
+ WL_TK_ACT[235] WL_TK_ACT[236] WL_TK_ACT[237] WL_TK_ACT[238] WL_TK_ACT[239] 
+ WL_TK_ACT[240] WL_TK_ACT[241] WL_TK_ACT[242] WL_TK_ACT[243] WL_TK_ACT[244] 
+ WL_TK_ACT[245] WL_TK_ACT[246] WL_TK_ACT[247] WL_TK_ACT[248] WL_TK_ACT[249] 
+ WL_TK_ACT[250] WL_TK_ACT[251] WL_TK_ACT[252] WL_TK_ACT[253] WL_TK_ACT[254] 
+ WL_TK_ACT[255] WL_TK_ACT[256] WL_TK_ACT[257] WL_TK_ACT[258] WL_TK_ACT[259] 
+ WL_TK_ACT[260] WL_TK_ACT[261] WL_TK_ACT[262] WL_TK_ACT[263] WL_TK_ACT[264] 
+ WL_TK_ACT[265] WL_TK_ACT[266] WL_TK_ACT[267] WL_TK_ACT[268] WL_TK_ACT[269] 
+ WL_TK_ACT[270] WL_TK_ACT[271] WL_TK_ACT[272] WL_TK_ACT[273] WL_TK_ACT[274] 
+ WL_TK_ACT[275] WL_TK_ACT[276] WL_TK_ACT[277] WL_TK_ACT[278] WL_TK_ACT[279] 
+ WL_TK_ACT[280] WL_TK_ACT[281] WL_TK_ACT[282] WL_TK_ACT[283] WL_TK_ACT[284] 
+ WL_TK_ACT[285] WL_TK_ACT[286] WL_TK_ACT[287] WL_TK_ACT[288] WL_TK_ACT[289] 
+ WL_TK_ACT[290] WL_TK_ACT[291] WL_TK_ACT[292] WL_TK_ACT[293] WL_TK_ACT[294] 
+ WL_TK_ACT[295] WL_TK_ACT[296] WL_TK_ACT[297] WL_TK_ACT[298] WL_TK_ACT[299] 
+ WL_TK_ACT[300] WL_TK_ACT[301] WL_TK_ACT[302] WL_TK_ACT[303] WL_TK_ACT[304] 
+ WL_TK_ACT[305] WL_TK_ACT[306] WL_TK_ACT[307] WL_TK_ACT[308] WL_TK_ACT[309] 
+ WL_TK_ACT[310] WL_TK_ACT[311] WL_TK_ACT[312] WL_TK_ACT[313] WL_TK_ACT[314] 
+ WL_TK_ACT[315] WL_TK_ACT[316] WL_TK_ACT[317] WL_TK_ACT[318] WL_TK_ACT[319] 
+ WL_TK_ACT[320] WL_TK_ACT[321] WL_TK_ACT[322] WL_TK_ACT[323] WL_TK_ACT[324] 
+ WL_TK_ACT[325] WL_TK_ACT[326] WL_TK_ACT[327] WL_TK_ACT[328] WL_TK_ACT[329] 
+ WL_TK_ACT[330] WL_TK_ACT[331] WL_TK_ACT[332] WL_TK_ACT[333] WL_TK_ACT[334] 
+ WL_TK_ACT[335] WL_TK_ACT[336] WL_TK_ACT[337] WL_TK_ACT[338] WL_TK_ACT[339] 
+ WL_TK_ACT[340] WL_TK_ACT[341] WL_TK_ACT[342] WL_TK_ACT[343] WL_TK_ACT[344] 
+ WL_TK_ACT[345] WL_TK_ACT[346] WL_TK_ACT[347] WL_TK_ACT[348] WL_TK_ACT[349] 
+ WL_TK_ACT[350] WL_TK_ACT[351] WL_TK_ACT[352] WL_TK_ACT[353] WL_TK_ACT[354] 
+ WL_TK_ACT[355] WL_TK_ACT[356] WL_TK_ACT[357] WL_TK_ACT[358] WL_TK_ACT[359] 
+ WL_TK_ACT[360] WL_TK_ACT[361] WL_TK_ACT[362] WL_TK_ACT[363] WL_TK_ACT[364] 
+ WL_TK_ACT[365] WL_TK_ACT[366] WL_TK_ACT[367] WL_TK_ACT[368] WL_TK_ACT[369] 
+ WL_TK_ACT[370] WL_TK_ACT[371] WL_TK_ACT[372] WL_TK_ACT[373] WL_TK_ACT[374] 
+ WL_TK_ACT[375] WL_TK_ACT[376] WL_TK_ACT[377] WL_TK_ACT[378] WL_TK_ACT[379] 
+ WL_TK_ACT[380] WL_TK_ACT[381] WL_TK_ACT[382] WL_TK_ACT[383] WL_TK_ACT[384] 
+ WL_TK_ACT[385] WL_TK_ACT[386] WL_TK_ACT[387] WL_TK_ACT[388] WL_TK_ACT[389] 
+ WL_TK_ACT[390] WL_TK_ACT[391] WL_TK_ACT[392] WL_TK_ACT[393] WL_TK_ACT[394] 
+ WL_TK_ACT[395] WL_TK_ACT[396] WL_TK_ACT[397] WL_TK_ACT[398] WL_TK_ACT[399] 
+ WL_TK_ACT[400] WL_TK_ACT[401] WL_TK_ACT[402] WL_TK_ACT[403] WL_TK_ACT[404] 
+ WL_TK_ACT[405] WL_TK_ACT[406] WL_TK_ACT[407] WL_TK_ACT[408] WL_TK_ACT[409] 
+ WL_TK_ACT[410] WL_TK_ACT[411] WL_TK_ACT[412] WL_TK_ACT[413] WL_TK_ACT[414] 
+ WL_TK_ACT[415] WL_TK_ACT[416] WL_TK_ACT[417] WL_TK_ACT[418] WL_TK_ACT[419] 
+ WL_TK_ACT[420] WL_TK_ACT[421] WL_TK_ACT[422] WL_TK_ACT[423] WL_TK_ACT[424] 
+ WL_TK_ACT[425] WL_TK_ACT[426] WL_TK_ACT[427] WL_TK_ACT[428] WL_TK_ACT[429] 
+ WL_TK_ACT[430] WL_TK_ACT[431] WL_TK_ACT[432] WL_TK_ACT[433] WL_TK_ACT[434] 
+ WL_TK_ACT[435] WL_TK_ACT[436] WL_TK_ACT[437] WL_TK_ACT[438] WL_TK_ACT[439] 
+ WL_TK_ACT[440] WL_TK_ACT[441] WL_TK_ACT[442] WL_TK_ACT[443] WL_TK_ACT[444] 
+ WL_TK_ACT[445] WL_TK_ACT[446] WL_TK_ACT[447] WL_TK_ACT[448] WL_TK_ACT[449] 
+ WL_TK_ACT[450] WL_TK_ACT[451] WL_TK_ACT[452] WL_TK_ACT[453] WL_TK_ACT[454] 
+ WL_TK_ACT[455] WL_TK_ACT[456] WL_TK_ACT[457] WL_TK_ACT[458] WL_TK_ACT[459] 
+ WL_TK_ACT[460] WL_TK_ACT[461] WL_TK_ACT[462] WL_TK_ACT[463] WL_TK_ACT[464] 
+ WL_TK_ACT[465] WL_TK_ACT[466] WL_TK_ACT[467] WL_TK_ACT[468] WL_TK_ACT[469] 
+ WL_TK_ACT[470] WL_TK_ACT[471] WL_TK_ACT[472] WL_TK_ACT[473] WL_TK_ACT[474] 
+ WL_TK_ACT[475] WL_TK_ACT[476] WL_TK_ACT[477] WL_TK_ACT[478] WL_TK_ACT[479] 
+ WL_TK_ACT[480] WL_TK_ACT[481] WL_TK_ACT[482] WL_TK_ACT[483] WL_TK_ACT[484] 
+ WL_TK_ACT[485] WL_TK_ACT[486] WL_TK_ACT[487] WL_TK_ACT[488] WL_TK_ACT[489] 
+ WL_TK_ACT[490] WL_TK_ACT[491] WL_TK_ACT[492] WL_TK_ACT[493] WL_TK_ACT[494] 
+ WL_TK_ACT[495] WL_TK_ACT[496] WL_TK_ACT[497] WL_TK_ACT[498] WL_TK_ACT[499] 
+ WL_TK_ACT[500] WL_TK_ACT[501] WL_TK_ACT[502] WL_TK_ACT[503] WL_TK_ACT[504] 
+ WL_TK_ACT[505] WL_TK_ACT[506] WL_TK_ACT[507] WL_TK_ACT[508] WL_TK_ACT[509] 
+ WL_TK_ACT[510] WL_TK_ACT[511] WL_TK_LD WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] 
+ X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] 
+ XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I BWEBM_LL:I BWEBM_LR:I BWEB_LL:I BWEB_LR:I CEB:I CEBM:I 
*.PININFO CLK:I DM_LL:I DM_LR:I D_LL:I D_LR:I PD:I PTSEL:I RTSEL[0]:I 
*.PININFO RTSEL[1]:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I 
*.PININFO X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I XM[0]:I 
*.PININFO XM[1]:I XM[2]:I XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I 
*.PININFO Y[0]:I Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I Q_LL:O 
*.PININFO Q_LR:O VDDI:B VSSI:B WL_TK_ACT[0]:B WL_TK_ACT[1]:B WL_TK_ACT[2]:B 
*.PININFO WL_TK_ACT[3]:B WL_TK_ACT[4]:B WL_TK_ACT[5]:B WL_TK_ACT[6]:B 
*.PININFO WL_TK_ACT[7]:B WL_TK_ACT[8]:B WL_TK_ACT[9]:B WL_TK_ACT[10]:B 
*.PININFO WL_TK_ACT[11]:B WL_TK_ACT[12]:B WL_TK_ACT[13]:B WL_TK_ACT[14]:B 
*.PININFO WL_TK_ACT[15]:B WL_TK_ACT[16]:B WL_TK_ACT[17]:B WL_TK_ACT[18]:B 
*.PININFO WL_TK_ACT[19]:B WL_TK_ACT[20]:B WL_TK_ACT[21]:B WL_TK_ACT[22]:B 
*.PININFO WL_TK_ACT[23]:B WL_TK_ACT[24]:B WL_TK_ACT[25]:B WL_TK_ACT[26]:B 
*.PININFO WL_TK_ACT[27]:B WL_TK_ACT[28]:B WL_TK_ACT[29]:B WL_TK_ACT[30]:B 
*.PININFO WL_TK_ACT[31]:B WL_TK_ACT[32]:B WL_TK_ACT[33]:B WL_TK_ACT[34]:B 
*.PININFO WL_TK_ACT[35]:B WL_TK_ACT[36]:B WL_TK_ACT[37]:B WL_TK_ACT[38]:B 
*.PININFO WL_TK_ACT[39]:B WL_TK_ACT[40]:B WL_TK_ACT[41]:B WL_TK_ACT[42]:B 
*.PININFO WL_TK_ACT[43]:B WL_TK_ACT[44]:B WL_TK_ACT[45]:B WL_TK_ACT[46]:B 
*.PININFO WL_TK_ACT[47]:B WL_TK_ACT[48]:B WL_TK_ACT[49]:B WL_TK_ACT[50]:B 
*.PININFO WL_TK_ACT[51]:B WL_TK_ACT[52]:B WL_TK_ACT[53]:B WL_TK_ACT[54]:B 
*.PININFO WL_TK_ACT[55]:B WL_TK_ACT[56]:B WL_TK_ACT[57]:B WL_TK_ACT[58]:B 
*.PININFO WL_TK_ACT[59]:B WL_TK_ACT[60]:B WL_TK_ACT[61]:B WL_TK_ACT[62]:B 
*.PININFO WL_TK_ACT[63]:B WL_TK_ACT[64]:B WL_TK_ACT[65]:B WL_TK_ACT[66]:B 
*.PININFO WL_TK_ACT[67]:B WL_TK_ACT[68]:B WL_TK_ACT[69]:B WL_TK_ACT[70]:B 
*.PININFO WL_TK_ACT[71]:B WL_TK_ACT[72]:B WL_TK_ACT[73]:B WL_TK_ACT[74]:B 
*.PININFO WL_TK_ACT[75]:B WL_TK_ACT[76]:B WL_TK_ACT[77]:B WL_TK_ACT[78]:B 
*.PININFO WL_TK_ACT[79]:B WL_TK_ACT[80]:B WL_TK_ACT[81]:B WL_TK_ACT[82]:B 
*.PININFO WL_TK_ACT[83]:B WL_TK_ACT[84]:B WL_TK_ACT[85]:B WL_TK_ACT[86]:B 
*.PININFO WL_TK_ACT[87]:B WL_TK_ACT[88]:B WL_TK_ACT[89]:B WL_TK_ACT[90]:B 
*.PININFO WL_TK_ACT[91]:B WL_TK_ACT[92]:B WL_TK_ACT[93]:B WL_TK_ACT[94]:B 
*.PININFO WL_TK_ACT[95]:B WL_TK_ACT[96]:B WL_TK_ACT[97]:B WL_TK_ACT[98]:B 
*.PININFO WL_TK_ACT[99]:B WL_TK_ACT[100]:B WL_TK_ACT[101]:B WL_TK_ACT[102]:B 
*.PININFO WL_TK_ACT[103]:B WL_TK_ACT[104]:B WL_TK_ACT[105]:B WL_TK_ACT[106]:B 
*.PININFO WL_TK_ACT[107]:B WL_TK_ACT[108]:B WL_TK_ACT[109]:B WL_TK_ACT[110]:B 
*.PININFO WL_TK_ACT[111]:B WL_TK_ACT[112]:B WL_TK_ACT[113]:B WL_TK_ACT[114]:B 
*.PININFO WL_TK_ACT[115]:B WL_TK_ACT[116]:B WL_TK_ACT[117]:B WL_TK_ACT[118]:B 
*.PININFO WL_TK_ACT[119]:B WL_TK_ACT[120]:B WL_TK_ACT[121]:B WL_TK_ACT[122]:B 
*.PININFO WL_TK_ACT[123]:B WL_TK_ACT[124]:B WL_TK_ACT[125]:B WL_TK_ACT[126]:B 
*.PININFO WL_TK_ACT[127]:B WL_TK_ACT[128]:B WL_TK_ACT[129]:B WL_TK_ACT[130]:B 
*.PININFO WL_TK_ACT[131]:B WL_TK_ACT[132]:B WL_TK_ACT[133]:B WL_TK_ACT[134]:B 
*.PININFO WL_TK_ACT[135]:B WL_TK_ACT[136]:B WL_TK_ACT[137]:B WL_TK_ACT[138]:B 
*.PININFO WL_TK_ACT[139]:B WL_TK_ACT[140]:B WL_TK_ACT[141]:B WL_TK_ACT[142]:B 
*.PININFO WL_TK_ACT[143]:B WL_TK_ACT[144]:B WL_TK_ACT[145]:B WL_TK_ACT[146]:B 
*.PININFO WL_TK_ACT[147]:B WL_TK_ACT[148]:B WL_TK_ACT[149]:B WL_TK_ACT[150]:B 
*.PININFO WL_TK_ACT[151]:B WL_TK_ACT[152]:B WL_TK_ACT[153]:B WL_TK_ACT[154]:B 
*.PININFO WL_TK_ACT[155]:B WL_TK_ACT[156]:B WL_TK_ACT[157]:B WL_TK_ACT[158]:B 
*.PININFO WL_TK_ACT[159]:B WL_TK_ACT[160]:B WL_TK_ACT[161]:B WL_TK_ACT[162]:B 
*.PININFO WL_TK_ACT[163]:B WL_TK_ACT[164]:B WL_TK_ACT[165]:B WL_TK_ACT[166]:B 
*.PININFO WL_TK_ACT[167]:B WL_TK_ACT[168]:B WL_TK_ACT[169]:B WL_TK_ACT[170]:B 
*.PININFO WL_TK_ACT[171]:B WL_TK_ACT[172]:B WL_TK_ACT[173]:B WL_TK_ACT[174]:B 
*.PININFO WL_TK_ACT[175]:B WL_TK_ACT[176]:B WL_TK_ACT[177]:B WL_TK_ACT[178]:B 
*.PININFO WL_TK_ACT[179]:B WL_TK_ACT[180]:B WL_TK_ACT[181]:B WL_TK_ACT[182]:B 
*.PININFO WL_TK_ACT[183]:B WL_TK_ACT[184]:B WL_TK_ACT[185]:B WL_TK_ACT[186]:B 
*.PININFO WL_TK_ACT[187]:B WL_TK_ACT[188]:B WL_TK_ACT[189]:B WL_TK_ACT[190]:B 
*.PININFO WL_TK_ACT[191]:B WL_TK_ACT[192]:B WL_TK_ACT[193]:B WL_TK_ACT[194]:B 
*.PININFO WL_TK_ACT[195]:B WL_TK_ACT[196]:B WL_TK_ACT[197]:B WL_TK_ACT[198]:B 
*.PININFO WL_TK_ACT[199]:B WL_TK_ACT[200]:B WL_TK_ACT[201]:B WL_TK_ACT[202]:B 
*.PININFO WL_TK_ACT[203]:B WL_TK_ACT[204]:B WL_TK_ACT[205]:B WL_TK_ACT[206]:B 
*.PININFO WL_TK_ACT[207]:B WL_TK_ACT[208]:B WL_TK_ACT[209]:B WL_TK_ACT[210]:B 
*.PININFO WL_TK_ACT[211]:B WL_TK_ACT[212]:B WL_TK_ACT[213]:B WL_TK_ACT[214]:B 
*.PININFO WL_TK_ACT[215]:B WL_TK_ACT[216]:B WL_TK_ACT[217]:B WL_TK_ACT[218]:B 
*.PININFO WL_TK_ACT[219]:B WL_TK_ACT[220]:B WL_TK_ACT[221]:B WL_TK_ACT[222]:B 
*.PININFO WL_TK_ACT[223]:B WL_TK_ACT[224]:B WL_TK_ACT[225]:B WL_TK_ACT[226]:B 
*.PININFO WL_TK_ACT[227]:B WL_TK_ACT[228]:B WL_TK_ACT[229]:B WL_TK_ACT[230]:B 
*.PININFO WL_TK_ACT[231]:B WL_TK_ACT[232]:B WL_TK_ACT[233]:B WL_TK_ACT[234]:B 
*.PININFO WL_TK_ACT[235]:B WL_TK_ACT[236]:B WL_TK_ACT[237]:B WL_TK_ACT[238]:B 
*.PININFO WL_TK_ACT[239]:B WL_TK_ACT[240]:B WL_TK_ACT[241]:B WL_TK_ACT[242]:B 
*.PININFO WL_TK_ACT[243]:B WL_TK_ACT[244]:B WL_TK_ACT[245]:B WL_TK_ACT[246]:B 
*.PININFO WL_TK_ACT[247]:B WL_TK_ACT[248]:B WL_TK_ACT[249]:B WL_TK_ACT[250]:B 
*.PININFO WL_TK_ACT[251]:B WL_TK_ACT[252]:B WL_TK_ACT[253]:B WL_TK_ACT[254]:B 
*.PININFO WL_TK_ACT[255]:B WL_TK_ACT[256]:B WL_TK_ACT[257]:B WL_TK_ACT[258]:B 
*.PININFO WL_TK_ACT[259]:B WL_TK_ACT[260]:B WL_TK_ACT[261]:B WL_TK_ACT[262]:B 
*.PININFO WL_TK_ACT[263]:B WL_TK_ACT[264]:B WL_TK_ACT[265]:B WL_TK_ACT[266]:B 
*.PININFO WL_TK_ACT[267]:B WL_TK_ACT[268]:B WL_TK_ACT[269]:B WL_TK_ACT[270]:B 
*.PININFO WL_TK_ACT[271]:B WL_TK_ACT[272]:B WL_TK_ACT[273]:B WL_TK_ACT[274]:B 
*.PININFO WL_TK_ACT[275]:B WL_TK_ACT[276]:B WL_TK_ACT[277]:B WL_TK_ACT[278]:B 
*.PININFO WL_TK_ACT[279]:B WL_TK_ACT[280]:B WL_TK_ACT[281]:B WL_TK_ACT[282]:B 
*.PININFO WL_TK_ACT[283]:B WL_TK_ACT[284]:B WL_TK_ACT[285]:B WL_TK_ACT[286]:B 
*.PININFO WL_TK_ACT[287]:B WL_TK_ACT[288]:B WL_TK_ACT[289]:B WL_TK_ACT[290]:B 
*.PININFO WL_TK_ACT[291]:B WL_TK_ACT[292]:B WL_TK_ACT[293]:B WL_TK_ACT[294]:B 
*.PININFO WL_TK_ACT[295]:B WL_TK_ACT[296]:B WL_TK_ACT[297]:B WL_TK_ACT[298]:B 
*.PININFO WL_TK_ACT[299]:B WL_TK_ACT[300]:B WL_TK_ACT[301]:B WL_TK_ACT[302]:B 
*.PININFO WL_TK_ACT[303]:B WL_TK_ACT[304]:B WL_TK_ACT[305]:B WL_TK_ACT[306]:B 
*.PININFO WL_TK_ACT[307]:B WL_TK_ACT[308]:B WL_TK_ACT[309]:B WL_TK_ACT[310]:B 
*.PININFO WL_TK_ACT[311]:B WL_TK_ACT[312]:B WL_TK_ACT[313]:B WL_TK_ACT[314]:B 
*.PININFO WL_TK_ACT[315]:B WL_TK_ACT[316]:B WL_TK_ACT[317]:B WL_TK_ACT[318]:B 
*.PININFO WL_TK_ACT[319]:B WL_TK_ACT[320]:B WL_TK_ACT[321]:B WL_TK_ACT[322]:B 
*.PININFO WL_TK_ACT[323]:B WL_TK_ACT[324]:B WL_TK_ACT[325]:B WL_TK_ACT[326]:B 
*.PININFO WL_TK_ACT[327]:B WL_TK_ACT[328]:B WL_TK_ACT[329]:B WL_TK_ACT[330]:B 
*.PININFO WL_TK_ACT[331]:B WL_TK_ACT[332]:B WL_TK_ACT[333]:B WL_TK_ACT[334]:B 
*.PININFO WL_TK_ACT[335]:B WL_TK_ACT[336]:B WL_TK_ACT[337]:B WL_TK_ACT[338]:B 
*.PININFO WL_TK_ACT[339]:B WL_TK_ACT[340]:B WL_TK_ACT[341]:B WL_TK_ACT[342]:B 
*.PININFO WL_TK_ACT[343]:B WL_TK_ACT[344]:B WL_TK_ACT[345]:B WL_TK_ACT[346]:B 
*.PININFO WL_TK_ACT[347]:B WL_TK_ACT[348]:B WL_TK_ACT[349]:B WL_TK_ACT[350]:B 
*.PININFO WL_TK_ACT[351]:B WL_TK_ACT[352]:B WL_TK_ACT[353]:B WL_TK_ACT[354]:B 
*.PININFO WL_TK_ACT[355]:B WL_TK_ACT[356]:B WL_TK_ACT[357]:B WL_TK_ACT[358]:B 
*.PININFO WL_TK_ACT[359]:B WL_TK_ACT[360]:B WL_TK_ACT[361]:B WL_TK_ACT[362]:B 
*.PININFO WL_TK_ACT[363]:B WL_TK_ACT[364]:B WL_TK_ACT[365]:B WL_TK_ACT[366]:B 
*.PININFO WL_TK_ACT[367]:B WL_TK_ACT[368]:B WL_TK_ACT[369]:B WL_TK_ACT[370]:B 
*.PININFO WL_TK_ACT[371]:B WL_TK_ACT[372]:B WL_TK_ACT[373]:B WL_TK_ACT[374]:B 
*.PININFO WL_TK_ACT[375]:B WL_TK_ACT[376]:B WL_TK_ACT[377]:B WL_TK_ACT[378]:B 
*.PININFO WL_TK_ACT[379]:B WL_TK_ACT[380]:B WL_TK_ACT[381]:B WL_TK_ACT[382]:B 
*.PININFO WL_TK_ACT[383]:B WL_TK_ACT[384]:B WL_TK_ACT[385]:B WL_TK_ACT[386]:B 
*.PININFO WL_TK_ACT[387]:B WL_TK_ACT[388]:B WL_TK_ACT[389]:B WL_TK_ACT[390]:B 
*.PININFO WL_TK_ACT[391]:B WL_TK_ACT[392]:B WL_TK_ACT[393]:B WL_TK_ACT[394]:B 
*.PININFO WL_TK_ACT[395]:B WL_TK_ACT[396]:B WL_TK_ACT[397]:B WL_TK_ACT[398]:B 
*.PININFO WL_TK_ACT[399]:B WL_TK_ACT[400]:B WL_TK_ACT[401]:B WL_TK_ACT[402]:B 
*.PININFO WL_TK_ACT[403]:B WL_TK_ACT[404]:B WL_TK_ACT[405]:B WL_TK_ACT[406]:B 
*.PININFO WL_TK_ACT[407]:B WL_TK_ACT[408]:B WL_TK_ACT[409]:B WL_TK_ACT[410]:B 
*.PININFO WL_TK_ACT[411]:B WL_TK_ACT[412]:B WL_TK_ACT[413]:B WL_TK_ACT[414]:B 
*.PININFO WL_TK_ACT[415]:B WL_TK_ACT[416]:B WL_TK_ACT[417]:B WL_TK_ACT[418]:B 
*.PININFO WL_TK_ACT[419]:B WL_TK_ACT[420]:B WL_TK_ACT[421]:B WL_TK_ACT[422]:B 
*.PININFO WL_TK_ACT[423]:B WL_TK_ACT[424]:B WL_TK_ACT[425]:B WL_TK_ACT[426]:B 
*.PININFO WL_TK_ACT[427]:B WL_TK_ACT[428]:B WL_TK_ACT[429]:B WL_TK_ACT[430]:B 
*.PININFO WL_TK_ACT[431]:B WL_TK_ACT[432]:B WL_TK_ACT[433]:B WL_TK_ACT[434]:B 
*.PININFO WL_TK_ACT[435]:B WL_TK_ACT[436]:B WL_TK_ACT[437]:B WL_TK_ACT[438]:B 
*.PININFO WL_TK_ACT[439]:B WL_TK_ACT[440]:B WL_TK_ACT[441]:B WL_TK_ACT[442]:B 
*.PININFO WL_TK_ACT[443]:B WL_TK_ACT[444]:B WL_TK_ACT[445]:B WL_TK_ACT[446]:B 
*.PININFO WL_TK_ACT[447]:B WL_TK_ACT[448]:B WL_TK_ACT[449]:B WL_TK_ACT[450]:B 
*.PININFO WL_TK_ACT[451]:B WL_TK_ACT[452]:B WL_TK_ACT[453]:B WL_TK_ACT[454]:B 
*.PININFO WL_TK_ACT[455]:B WL_TK_ACT[456]:B WL_TK_ACT[457]:B WL_TK_ACT[458]:B 
*.PININFO WL_TK_ACT[459]:B WL_TK_ACT[460]:B WL_TK_ACT[461]:B WL_TK_ACT[462]:B 
*.PININFO WL_TK_ACT[463]:B WL_TK_ACT[464]:B WL_TK_ACT[465]:B WL_TK_ACT[466]:B 
*.PININFO WL_TK_ACT[467]:B WL_TK_ACT[468]:B WL_TK_ACT[469]:B WL_TK_ACT[470]:B 
*.PININFO WL_TK_ACT[471]:B WL_TK_ACT[472]:B WL_TK_ACT[473]:B WL_TK_ACT[474]:B 
*.PININFO WL_TK_ACT[475]:B WL_TK_ACT[476]:B WL_TK_ACT[477]:B WL_TK_ACT[478]:B 
*.PININFO WL_TK_ACT[479]:B WL_TK_ACT[480]:B WL_TK_ACT[481]:B WL_TK_ACT[482]:B 
*.PININFO WL_TK_ACT[483]:B WL_TK_ACT[484]:B WL_TK_ACT[485]:B WL_TK_ACT[486]:B 
*.PININFO WL_TK_ACT[487]:B WL_TK_ACT[488]:B WL_TK_ACT[489]:B WL_TK_ACT[490]:B 
*.PININFO WL_TK_ACT[491]:B WL_TK_ACT[492]:B WL_TK_ACT[493]:B WL_TK_ACT[494]:B 
*.PININFO WL_TK_ACT[495]:B WL_TK_ACT[496]:B WL_TK_ACT[497]:B WL_TK_ACT[498]:B 
*.PININFO WL_TK_ACT[499]:B WL_TK_ACT[500]:B WL_TK_ACT[501]:B WL_TK_ACT[502]:B 
*.PININFO WL_TK_ACT[503]:B WL_TK_ACT[504]:B WL_TK_ACT[505]:B WL_TK_ACT[506]:B 
*.PININFO WL_TK_ACT[507]:B WL_TK_ACT[508]:B WL_TK_ACT[509]:B WL_TK_ACT[510]:B 
*.PININFO WL_TK_ACT[511]:B WL_TK_LD:B
XARR_WLLD_RD VDDI VDDHD VDDI VSSI WL_RD2[0] WL_RD2[1] WL_RD3[0] WL_RD3[1] 
+ S1AHSF400W40_SB_ARR_WLLD_SIM
XARR_WLLD_RU VDDI VDDHD VDDI VSSI WL_RU2[0] WL_RU2[1] WL_RU3[0] WL_RU3[1] 
+ S1AHSF400W40_SB_ARR_WLLD_SIM
XARR_WLLD_LD VDDI VDDHD VDDI VSSI WL_LD3[0] WL_LD3[1] WL_LD2[0] WL_LD2[1] 
+ S1AHSF400W40_SB_ARR_WLLD_SIM
XARR_WLLD_LU VDDI VDDHD VDDI VSSI WL_LU3[0] WL_LU3[1] WL_LU2[0] WL_LU2[1] 
+ S1AHSF400W40_SB_ARR_WLLD_SIM
XARR_BLLD_LL BLB_LL_2 BLB_LL_3 BL_LL_2 BL_LL_3 VDDI VSSI S1AHSF400W40_SB_ARR_BLLD_SIM
XARR_BLLD_LR BLB_LR_2 BLB_LR_3 BL_LR_2 BL_LR_3 VDDI VSSI S1AHSF400W40_SB_ARR_BLLD_SIM
XBK_STRAP_U DEC_X0_21[0] DEC_X0_21[1] DEC_X0_21[2] DEC_X0_21[3] DEC_X0_21[4] 
+ DEC_X0_21[5] DEC_X0_21[6] DEC_X0_21[7] DEC_X0_22[0] DEC_X0_22[1] 
+ DEC_X0_22[2] DEC_X0_22[3] DEC_X0_22[4] DEC_X0_22[5] DEC_X0_22[6] 
+ DEC_X0_22[7] DEC_X1_21[0] DEC_X1_21[1] DEC_X1_21[2] DEC_X1_21[3] 
+ DEC_X1_21[4] DEC_X1_21[5] DEC_X1_21[6] DEC_X1_21[7] DEC_X1_22[0] 
+ DEC_X1_22[1] DEC_X1_22[2] DEC_X1_22[3] DEC_X1_22[4] DEC_X1_22[5] 
+ DEC_X1_22[6] DEC_X1_22[7] DEC_X2_21[0] DEC_X2_21[1] DEC_X2_21[2] 
+ DEC_X2_21[3] DEC_X2_21[4] DEC_X2_21[5] DEC_X2_21[6] DEC_X2_21[7] 
+ DEC_X2_SHARE_22 DEC_X2_22[0] DEC_X2_22[1] DEC_X2_22[2] DEC_X2_22[3] 
+ DEC_X2_22[4] DEC_X2_22[5] DEC_X2_22[6] DEC_X2_22[7] PD_BUF_21 PD_BUF_22 
+ VDDHD VDDI VSSI S1AHSF400W40_SB_STRAP_U_SIM
XTKBL TRKBL BL_TK_TP VDDHD PD VDDHD VDDI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI WL_TK_ACT[0] 
+ WL_TK_ACT[1] WL_TK_ACT[2] WL_TK_ACT[3] WL_TK_ACT[4] WL_TK_ACT[5] 
+ WL_TK_ACT[6] WL_TK_ACT[7] WL_TK_ACT[8] WL_TK_ACT[9] WL_TK_ACT[10] 
+ WL_TK_ACT[11] WL_TK_ACT[12] WL_TK_ACT[13] WL_TK_ACT[14] WL_TK_ACT[15] 
+ WL_TK_ACT[16] WL_TK_ACT[17] WL_TK_ACT[18] WL_TK_ACT[19] WL_TK_ACT[20] 
+ WL_TK_ACT[21] WL_TK_ACT[22] WL_TK_ACT[23] WL_TK_ACT[24] WL_TK_ACT[25] 
+ WL_TK_ACT[26] WL_TK_ACT[27] WL_TK_ACT[28] WL_TK_ACT[29] WL_TK_ACT[30] 
+ WL_TK_ACT[31] WL_TK_ACT[32] WL_TK_ACT[33] WL_TK_ACT[34] WL_TK_ACT[35] 
+ WL_TK_ACT[36] WL_TK_ACT[37] WL_TK_ACT[38] WL_TK_ACT[39] WL_TK_ACT[40] 
+ WL_TK_ACT[41] WL_TK_ACT[42] WL_TK_ACT[43] WL_TK_ACT[44] WL_TK_ACT[45] 
+ WL_TK_ACT[46] WL_TK_ACT[47] WL_TK_ACT[48] WL_TK_ACT[49] WL_TK_ACT[50] 
+ WL_TK_ACT[51] WL_TK_ACT[52] WL_TK_ACT[53] WL_TK_ACT[54] WL_TK_ACT[55] 
+ WL_TK_ACT[56] WL_TK_ACT[57] WL_TK_ACT[58] WL_TK_ACT[59] WL_TK_ACT[60] 
+ WL_TK_ACT[61] WL_TK_ACT[62] WL_TK_ACT[63] WL_TK_ACT[64] WL_TK_ACT[65] 
+ WL_TK_ACT[66] WL_TK_ACT[67] WL_TK_ACT[68] WL_TK_ACT[69] WL_TK_ACT[70] 
+ WL_TK_ACT[71] WL_TK_ACT[72] WL_TK_ACT[73] WL_TK_ACT[74] WL_TK_ACT[75] 
+ WL_TK_ACT[76] WL_TK_ACT[77] WL_TK_ACT[78] WL_TK_ACT[79] WL_TK_ACT[80] 
+ WL_TK_ACT[81] WL_TK_ACT[82] WL_TK_ACT[83] WL_TK_ACT[84] WL_TK_ACT[85] 
+ WL_TK_ACT[86] WL_TK_ACT[87] WL_TK_ACT[88] WL_TK_ACT[89] WL_TK_ACT[90] 
+ WL_TK_ACT[91] WL_TK_ACT[92] WL_TK_ACT[93] WL_TK_ACT[94] WL_TK_ACT[95] 
+ WL_TK_ACT[96] WL_TK_ACT[97] WL_TK_ACT[98] WL_TK_ACT[99] WL_TK_ACT[100] 
+ WL_TK_ACT[101] WL_TK_ACT[102] WL_TK_ACT[103] WL_TK_ACT[104] WL_TK_ACT[105] 
+ WL_TK_ACT[106] WL_TK_ACT[107] WL_TK_ACT[108] WL_TK_ACT[109] WL_TK_ACT[110] 
+ WL_TK_ACT[111] WL_TK_ACT[112] WL_TK_ACT[113] WL_TK_ACT[114] WL_TK_ACT[115] 
+ WL_TK_ACT[116] WL_TK_ACT[117] WL_TK_ACT[118] WL_TK_ACT[119] WL_TK_ACT[120] 
+ WL_TK_ACT[121] WL_TK_ACT[122] WL_TK_ACT[123] WL_TK_ACT[124] WL_TK_ACT[125] 
+ WL_TK_ACT[126] WL_TK_ACT[127] WL_TK_ACT[128] WL_TK_ACT[129] WL_TK_ACT[130] 
+ WL_TK_ACT[131] WL_TK_ACT[132] WL_TK_ACT[133] WL_TK_ACT[134] WL_TK_ACT[135] 
+ WL_TK_ACT[136] WL_TK_ACT[137] WL_TK_ACT[138] WL_TK_ACT[139] WL_TK_ACT[140] 
+ WL_TK_ACT[141] WL_TK_ACT[142] WL_TK_ACT[143] WL_TK_ACT[144] WL_TK_ACT[145] 
+ WL_TK_ACT[146] WL_TK_ACT[147] WL_TK_ACT[148] WL_TK_ACT[149] WL_TK_ACT[150] 
+ WL_TK_ACT[151] WL_TK_ACT[152] WL_TK_ACT[153] WL_TK_ACT[154] WL_TK_ACT[155] 
+ WL_TK_ACT[156] WL_TK_ACT[157] WL_TK_ACT[158] WL_TK_ACT[159] WL_TK_ACT[160] 
+ WL_TK_ACT[161] WL_TK_ACT[162] WL_TK_ACT[163] WL_TK_ACT[164] WL_TK_ACT[165] 
+ WL_TK_ACT[166] WL_TK_ACT[167] WL_TK_ACT[168] WL_TK_ACT[169] WL_TK_ACT[170] 
+ WL_TK_ACT[171] WL_TK_ACT[172] WL_TK_ACT[173] WL_TK_ACT[174] WL_TK_ACT[175] 
+ WL_TK_ACT[176] WL_TK_ACT[177] WL_TK_ACT[178] WL_TK_ACT[179] WL_TK_ACT[180] 
+ WL_TK_ACT[181] WL_TK_ACT[182] WL_TK_ACT[183] WL_TK_ACT[184] WL_TK_ACT[185] 
+ WL_TK_ACT[186] WL_TK_ACT[187] WL_TK_ACT[188] WL_TK_ACT[189] WL_TK_ACT[190] 
+ WL_TK_ACT[191] WL_TK_ACT[192] WL_TK_ACT[193] WL_TK_ACT[194] WL_TK_ACT[195] 
+ WL_TK_ACT[196] WL_TK_ACT[197] WL_TK_ACT[198] WL_TK_ACT[199] WL_TK_ACT[200] 
+ WL_TK_ACT[201] WL_TK_ACT[202] WL_TK_ACT[203] WL_TK_ACT[204] WL_TK_ACT[205] 
+ WL_TK_ACT[206] WL_TK_ACT[207] WL_TK_ACT[208] WL_TK_ACT[209] WL_TK_ACT[210] 
+ WL_TK_ACT[211] WL_TK_ACT[212] WL_TK_ACT[213] WL_TK_ACT[214] WL_TK_ACT[215] 
+ WL_TK_ACT[216] WL_TK_ACT[217] WL_TK_ACT[218] WL_TK_ACT[219] WL_TK_ACT[220] 
+ WL_TK_ACT[221] WL_TK_ACT[222] WL_TK_ACT[223] WL_TK_ACT[224] WL_TK_ACT[225] 
+ WL_TK_ACT[226] WL_TK_ACT[227] WL_TK_ACT[228] WL_TK_ACT[229] WL_TK_ACT[230] 
+ WL_TK_ACT[231] WL_TK_ACT[232] WL_TK_ACT[233] WL_TK_ACT[234] WL_TK_ACT[235] 
+ WL_TK_ACT[236] WL_TK_ACT[237] WL_TK_ACT[238] WL_TK_ACT[239] WL_TK_ACT[240] 
+ WL_TK_ACT[241] WL_TK_ACT[242] WL_TK_ACT[243] WL_TK_ACT[244] WL_TK_ACT[245] 
+ WL_TK_ACT[246] WL_TK_ACT[247] WL_TK_ACT[248] WL_TK_ACT[249] WL_TK_ACT[250] 
+ WL_TK_ACT[251] WL_TK_ACT[252] WL_TK_ACT[253] WL_TK_ACT[254] WL_TK_ACT[255] 
+ WL_TK_ACT[256] WL_TK_ACT[257] WL_TK_ACT[258] WL_TK_ACT[259] WL_TK_ACT[260] 
+ WL_TK_ACT[261] WL_TK_ACT[262] WL_TK_ACT[263] WL_TK_ACT[264] WL_TK_ACT[265] 
+ WL_TK_ACT[266] WL_TK_ACT[267] WL_TK_ACT[268] WL_TK_ACT[269] WL_TK_ACT[270] 
+ WL_TK_ACT[271] WL_TK_ACT[272] WL_TK_ACT[273] WL_TK_ACT[274] WL_TK_ACT[275] 
+ WL_TK_ACT[276] WL_TK_ACT[277] WL_TK_ACT[278] WL_TK_ACT[279] WL_TK_ACT[280] 
+ WL_TK_ACT[281] WL_TK_ACT[282] WL_TK_ACT[283] WL_TK_ACT[284] WL_TK_ACT[285] 
+ WL_TK_ACT[286] WL_TK_ACT[287] WL_TK_ACT[288] WL_TK_ACT[289] WL_TK_ACT[290] 
+ WL_TK_ACT[291] WL_TK_ACT[292] WL_TK_ACT[293] WL_TK_ACT[294] WL_TK_ACT[295] 
+ WL_TK_ACT[296] WL_TK_ACT[297] WL_TK_ACT[298] WL_TK_ACT[299] WL_TK_ACT[300] 
+ WL_TK_ACT[301] WL_TK_ACT[302] WL_TK_ACT[303] WL_TK_ACT[304] WL_TK_ACT[305] 
+ WL_TK_ACT[306] WL_TK_ACT[307] WL_TK_ACT[308] WL_TK_ACT[309] WL_TK_ACT[310] 
+ WL_TK_ACT[311] WL_TK_ACT[312] WL_TK_ACT[313] WL_TK_ACT[314] WL_TK_ACT[315] 
+ WL_TK_ACT[316] WL_TK_ACT[317] WL_TK_ACT[318] WL_TK_ACT[319] WL_TK_ACT[320] 
+ WL_TK_ACT[321] WL_TK_ACT[322] WL_TK_ACT[323] WL_TK_ACT[324] WL_TK_ACT[325] 
+ WL_TK_ACT[326] WL_TK_ACT[327] WL_TK_ACT[328] WL_TK_ACT[329] WL_TK_ACT[330] 
+ WL_TK_ACT[331] WL_TK_ACT[332] WL_TK_ACT[333] WL_TK_ACT[334] WL_TK_ACT[335] 
+ WL_TK_ACT[336] WL_TK_ACT[337] WL_TK_ACT[338] WL_TK_ACT[339] WL_TK_ACT[340] 
+ WL_TK_ACT[341] WL_TK_ACT[342] WL_TK_ACT[343] WL_TK_ACT[344] WL_TK_ACT[345] 
+ WL_TK_ACT[346] WL_TK_ACT[347] WL_TK_ACT[348] WL_TK_ACT[349] WL_TK_ACT[350] 
+ WL_TK_ACT[351] WL_TK_ACT[352] WL_TK_ACT[353] WL_TK_ACT[354] WL_TK_ACT[355] 
+ WL_TK_ACT[356] WL_TK_ACT[357] WL_TK_ACT[358] WL_TK_ACT[359] WL_TK_ACT[360] 
+ WL_TK_ACT[361] WL_TK_ACT[362] WL_TK_ACT[363] WL_TK_ACT[364] WL_TK_ACT[365] 
+ WL_TK_ACT[366] WL_TK_ACT[367] WL_TK_ACT[368] WL_TK_ACT[369] WL_TK_ACT[370] 
+ WL_TK_ACT[371] WL_TK_ACT[372] WL_TK_ACT[373] WL_TK_ACT[374] WL_TK_ACT[375] 
+ WL_TK_ACT[376] WL_TK_ACT[377] WL_TK_ACT[378] WL_TK_ACT[379] WL_TK_ACT[380] 
+ WL_TK_ACT[381] WL_TK_ACT[382] WL_TK_ACT[383] WL_TK_ACT[384] WL_TK_ACT[385] 
+ WL_TK_ACT[386] WL_TK_ACT[387] WL_TK_ACT[388] WL_TK_ACT[389] WL_TK_ACT[390] 
+ WL_TK_ACT[391] WL_TK_ACT[392] WL_TK_ACT[393] WL_TK_ACT[394] WL_TK_ACT[395] 
+ WL_TK_ACT[396] WL_TK_ACT[397] WL_TK_ACT[398] WL_TK_ACT[399] WL_TK_ACT[400] 
+ WL_TK_ACT[401] WL_TK_ACT[402] WL_TK_ACT[403] WL_TK_ACT[404] WL_TK_ACT[405] 
+ WL_TK_ACT[406] WL_TK_ACT[407] WL_TK_ACT[408] WL_TK_ACT[409] WL_TK_ACT[410] 
+ WL_TK_ACT[411] WL_TK_ACT[412] WL_TK_ACT[413] WL_TK_ACT[414] WL_TK_ACT[415] 
+ WL_TK_ACT[416] WL_TK_ACT[417] WL_TK_ACT[418] WL_TK_ACT[419] WL_TK_ACT[420] 
+ WL_TK_ACT[421] WL_TK_ACT[422] WL_TK_ACT[423] WL_TK_ACT[424] WL_TK_ACT[425] 
+ WL_TK_ACT[426] WL_TK_ACT[427] WL_TK_ACT[428] WL_TK_ACT[429] WL_TK_ACT[430] 
+ WL_TK_ACT[431] WL_TK_ACT[432] WL_TK_ACT[433] WL_TK_ACT[434] WL_TK_ACT[435] 
+ WL_TK_ACT[436] WL_TK_ACT[437] WL_TK_ACT[438] WL_TK_ACT[439] WL_TK_ACT[440] 
+ WL_TK_ACT[441] WL_TK_ACT[442] WL_TK_ACT[443] WL_TK_ACT[444] WL_TK_ACT[445] 
+ WL_TK_ACT[446] WL_TK_ACT[447] WL_TK_ACT[448] WL_TK_ACT[449] WL_TK_ACT[450] 
+ WL_TK_ACT[451] WL_TK_ACT[452] WL_TK_ACT[453] WL_TK_ACT[454] WL_TK_ACT[455] 
+ WL_TK_ACT[456] WL_TK_ACT[457] WL_TK_ACT[458] WL_TK_ACT[459] WL_TK_ACT[460] 
+ WL_TK_ACT[461] WL_TK_ACT[462] WL_TK_ACT[463] WL_TK_ACT[464] WL_TK_ACT[465] 
+ WL_TK_ACT[466] WL_TK_ACT[467] WL_TK_ACT[468] WL_TK_ACT[469] WL_TK_ACT[470] 
+ WL_TK_ACT[471] WL_TK_ACT[472] WL_TK_ACT[473] WL_TK_ACT[474] WL_TK_ACT[475] 
+ WL_TK_ACT[476] WL_TK_ACT[477] WL_TK_ACT[478] WL_TK_ACT[479] WL_TK_ACT[480] 
+ WL_TK_ACT[481] WL_TK_ACT[482] WL_TK_ACT[483] WL_TK_ACT[484] WL_TK_ACT[485] 
+ WL_TK_ACT[486] WL_TK_ACT[487] WL_TK_ACT[488] WL_TK_ACT[489] WL_TK_ACT[490] 
+ WL_TK_ACT[491] WL_TK_ACT[492] WL_TK_ACT[493] WL_TK_ACT[494] WL_TK_ACT[495] 
+ WL_TK_ACT[496] WL_TK_ACT[497] WL_TK_ACT[498] WL_TK_ACT[499] WL_TK_ACT[500] 
+ WL_TK_ACT[501] WL_TK_ACT[502] WL_TK_ACT[503] WL_TK_ACT[504] WL_TK_ACT[505] 
+ WL_TK_ACT[506] WL_TK_ACT[507] WL_TK_ACT[508] WL_TK_ACT[509] WL_TK_ACT[510] 
+ WL_TK_ACT[511] TIEH_BT TIEL S1AHSF400W40_TKBL_SIM
XTRKPRE PD TRKBL WL_TK VDDHD VDDI VSSI TIEH_BT TIEL S1AHSF400W40_TRKPRE_SIM
XBK_WLDV_D DEC_X0_1[0] DEC_X0_1[1] DEC_X0_1[2] DEC_X0_1[3] DEC_X0_1[4] 
+ DEC_X0_1[5] DEC_X0_1[6] DEC_X0_1[7] DEC_X0_2[0] DEC_X0_2[1] DEC_X0_2[2] 
+ DEC_X0_2[3] DEC_X0_2[4] DEC_X0_2[5] DEC_X0_2[6] DEC_X0_2[7] DEC_X1_1[0] 
+ DEC_X1_1[1] DEC_X1_1[2] DEC_X1_1[3] DEC_X1_1[4] DEC_X1_1[5] DEC_X1_1[6] 
+ DEC_X1_1[7] DEC_X1_2[0] DEC_X1_2[1] DEC_X1_2[2] DEC_X1_2[3] DEC_X1_2[4] 
+ DEC_X1_2[5] DEC_X1_2[6] DEC_X1_2[7] DEC_X2_1[0] DEC_X2_1[1] DEC_X2_1[2] 
+ DEC_X2_1[3] DEC_X2_1[4] DEC_X2_1[5] DEC_X2_1[6] DEC_X2_1[7] DEC_X2_SHARE_2 
+ DEC_X2_2[0] DEC_X2_2[1] DEC_X2_2[2] DEC_X2_2[3] DEC_X2_2[4] DEC_X2_2[5] 
+ DEC_X2_2[6] DEC_X2_2[7] PD_BUF_L1 PD_BUF_2 VDDHD VDDI VSSI WL_LD1[0] 
+ WL_LD1[1] WL_RD1[0] WL_RD1[1] S1AHSF400W40_SB_WLDV_D_SIM
XBK_WLDV_U DEC_X0_3[0] DEC_X0_3[1] DEC_X0_3[2] DEC_X0_3[3] DEC_X0_3[4] 
+ DEC_X0_3[5] DEC_X0_3[6] DEC_X0_3[7] NET0528[0] NET0528[1] NET0528[2] 
+ NET0528[3] NET0528[4] NET0528[5] NET0528[6] NET0528[7] DEC_X1_3[0] 
+ DEC_X1_3[1] DEC_X1_3[2] DEC_X1_3[3] DEC_X1_3[4] DEC_X1_3[5] DEC_X1_3[6] 
+ DEC_X1_3[7] NET0527[0] NET0527[1] NET0527[2] NET0527[3] NET0527[4] 
+ NET0527[5] NET0527[6] NET0527[7] DEC_X2_3[0] DEC_X2_3[1] DEC_X2_3[2] 
+ DEC_X2_3[3] DEC_X2_3[4] DEC_X2_3[5] DEC_X2_3[6] DEC_X2_3[7] DEC_X2_SHARE_3 
+ NET0152 NET0525[0] NET0525[1] NET0525[2] NET0525[3] NET0525[4] NET0525[5] 
+ NET0525[6] NET0525[7] PD_BUF_3 NET0526 VDDHD VDDI VSSI WL_LU1[0] WL_LU1[1] 
+ WL_RU1[0] WL_RU1[1] S1AHSF400W40_SB_WLDV_U_SIM
XBK_WLDV_LD_U DEC_X0_22[0] DEC_X0_22[1] DEC_X0_22[2] DEC_X0_22[3] DEC_X0_22[4] 
+ DEC_X0_22[5] DEC_X0_22[6] DEC_X0_22[7] DEC_X0_3[0] DEC_X0_3[1] DEC_X0_3[2] 
+ DEC_X0_3[3] DEC_X0_3[4] DEC_X0_3[5] DEC_X0_3[6] DEC_X0_3[7] DEC_X1_22[0] 
+ DEC_X1_22[1] DEC_X1_22[2] DEC_X1_22[3] DEC_X1_22[4] DEC_X1_22[5] 
+ DEC_X1_22[6] DEC_X1_22[7] DEC_X1_3[0] DEC_X1_3[1] DEC_X1_3[2] DEC_X1_3[3] 
+ DEC_X1_3[4] DEC_X1_3[5] DEC_X1_3[6] DEC_X1_3[7] DEC_X2_22[0] DEC_X2_22[1] 
+ DEC_X2_22[2] DEC_X2_22[3] DEC_X2_22[4] DEC_X2_22[5] DEC_X2_22[6] 
+ DEC_X2_22[7] DEC_X2_SHARE_22 DEC_X2_SHARE_3 DEC_X2_3[0] DEC_X2_3[1] 
+ DEC_X2_3[2] DEC_X2_3[3] DEC_X2_3[4] DEC_X2_3[5] DEC_X2_3[6] DEC_X2_3[7] 
+ PD_BUF_22 PD_BUF_3 VDDHD VDDI VSSI S1AHSF400W40_SB_BK_LD_U_SIM
XARR_MCB_RDR NET142 NET143 NET144 NET141 VDDI VDDHD VDDI VSSI WL_RD3[0] 
+ WL_RD3[1] WL_RD4[0] WL_RD4[1] S1AHSF400W40_SB_ARR_MCB_SIM
XARR_MCB_LUR BLB_LR_3 NET0530 BL_LR_3 NET0190 VDDI VDDHD VDDI VSSI WL_LU2[0] 
+ WL_LU2[1] WL_LU1[0] WL_LU1[1] S1AHSF400W40_SB_ARR_MCB_SIM
XARR_MCB_RUL NET162 NET163 NET164 NET161 VDDI VDDHD VDDI VSSI WL_RU1[0] 
+ WL_RU1[1] WL_RU2[0] WL_RU2[1] S1AHSF400W40_SB_ARR_MCB_SIM
XARR_MCB_RUR NET172 NET173 NET174 NET565 VDDI VDDHD VDDI VSSI WL_RU3[0] 
+ WL_RU3[1] WL_RU4[0] WL_RU4[1] S1AHSF400W40_SB_ARR_MCB_SIM
XARR_MCB_RDL NET571 NET542 NET541 NET545 VDDI VDDHD VDDI VSSI WL_RD1[0] 
+ WL_RD1[1] WL_RD2[0] WL_RD2[1] S1AHSF400W40_SB_ARR_MCB_SIM
XARR_MCB_LDL BLB_LL_1[0] BLB_LL_2 BL_LL_1[0] BL_LL_2 VDDI VDDHD VDDI VSSI 
+ WL_LD4[0] WL_LD4[1] WL_LD3[0] WL_LD3[1] S1AHSF400W40_SB_ARR_MCB_SIM
XARR_MCB_LUL BLB_LL_3 NET0531 BL_LL_3 NET0240 VDDI VDDHD VDDI VSSI WL_LU4[0] 
+ WL_LU4[1] WL_LU3[0] WL_LU3[1] S1AHSF400W40_SB_ARR_MCB_SIM
XARR_MCB_LDR BLB_LR_1[0] BLB_LR_2 BL_LR_1[0] BL_LR_2 VDDI VDDHD VDDI VSSI 
+ WL_LD2[0] WL_LD2[1] WL_LD1[0] WL_LD1[1] S1AHSF400W40_SB_ARR_MCB_SIM
XBK_WLDV_LD_D DEC_X0_2[0] DEC_X0_2[1] DEC_X0_2[2] DEC_X0_2[3] DEC_X0_2[4] 
+ DEC_X0_2[5] DEC_X0_2[6] DEC_X0_2[7] DEC_X0_21[0] DEC_X0_21[1] DEC_X0_21[2] 
+ DEC_X0_21[3] DEC_X0_21[4] DEC_X0_21[5] DEC_X0_21[6] DEC_X0_21[7] DEC_X1_2[0] 
+ DEC_X1_2[1] DEC_X1_2[2] DEC_X1_2[3] DEC_X1_2[4] DEC_X1_2[5] DEC_X1_2[6] 
+ DEC_X1_2[7] DEC_X1_21[0] DEC_X1_21[1] DEC_X1_21[2] DEC_X1_21[3] DEC_X1_21[4] 
+ DEC_X1_21[5] DEC_X1_21[6] DEC_X1_21[7] DEC_X2_2[0] DEC_X2_2[1] DEC_X2_2[2] 
+ DEC_X2_2[3] DEC_X2_2[4] DEC_X2_2[5] DEC_X2_2[6] DEC_X2_2[7] DEC_X2_SHARE_2 
+ DEC_X2_21[0] DEC_X2_21[1] DEC_X2_21[2] DEC_X2_21[3] DEC_X2_21[4] 
+ DEC_X2_21[5] DEC_X2_21[6] DEC_X2_21[7] PD_BUF_2 PD_BUF_21 VDDHD VDDI VSSI 
+ S1AHSF400W40_SB_BK_LD_SIM
XIO_LD_L AWT2_L3 AWT2_L2 BIST2IO_L3 BIST2IO_L2 BLEQ_L3 BLEQ_L2 CKD_L3 CKD_L2 
+ PD_BUF_L3 PD_BUF_L2 RE_L3 RE_L2 SAE_L3 SAE_L2 VDDHD VDDI VSSI WE_L3 WE_L2 
+ YL_L3[0] YL_L3[1] YL_L2[0] YL_L2[1] DEC_Y_L3[0] DEC_Y_L3[1] DEC_Y_L3[2] 
+ DEC_Y_L3[3] DEC_Y_L3[4] DEC_Y_L3[5] DEC_Y_L3[6] DEC_Y_L3[7] DEC_Y_L2[0] 
+ DEC_Y_L2[1] DEC_Y_L2[2] DEC_Y_L2[3] DEC_Y_L2[4] DEC_Y_L2[5] DEC_Y_L2[6] 
+ DEC_Y_L2[7] S1AHSF400W40_SB_IO_LD_SIM
XIO_LD_R AWT2_R2 AWT2_R3 BIST2IO_R2 BIST2IO_R3 BLEQ_R2 BLEQ_R3 CKD_R2 CKD_R3 
+ PD_BUF_R2 PD_BUF_R3 RE_R2 RE_R3 SAE_R2 SAE_R3 VDDHD VDDI VSSI WE_R2 WE_R3 
+ YL_R2[0] YL_R2[1] YL_R3[0] YL_R3[1] DEC_Y_R2[0] DEC_Y_R2[1] DEC_Y_R2[2] 
+ DEC_Y_R2[3] DEC_Y_R2[4] DEC_Y_R2[5] DEC_Y_R2[6] DEC_Y_R2[7] DEC_Y_R3[0] 
+ DEC_Y_R3[1] DEC_Y_R3[2] DEC_Y_R3[3] DEC_Y_R3[4] DEC_Y_R3[5] DEC_Y_R3[6] 
+ DEC_Y_R3[7] S1AHSF400W40_SB_IO_LD_SIM
XIO_RR AWT2_R3 AWT2_R4 BIST2IO_R3 BIST2IO_R4 NET0545[0] NET0545[1] NET0545[2] 
+ NET0545[3] NET0545[4] NET0545[5] NET0545[6] NET0545[7] NET0545[8] NET0545[9] 
+ NET0545[10] NET0545[11] NET0545[12] NET0545[13] NET0545[14] NET0545[15] 
+ NET0544[0] NET0544[1] NET0544[2] NET0544[3] NET0544[4] NET0544[5] NET0544[6] 
+ NET0544[7] NET0544[8] NET0544[9] NET0544[10] NET0544[11] NET0544[12] 
+ NET0544[13] NET0544[14] NET0544[15] BLEQ_R3 BLEQ_R4 NET0543 NET0542 CKD_R3 
+ CKD_R4 NET0541 NET0540 PD_BUF_R3 PD_BUF_R4 NET0539 RE_R3 RE_R4 SAE_R3 SAE_R4 
+ VDDHD VDDI VSSI WE_R3 WE_R4 YL_R3[0] YL_R3[1] YL_R4[0] YL_R4[1] DEC_Y_R3[0] 
+ DEC_Y_R3[1] DEC_Y_R3[2] DEC_Y_R3[3] DEC_Y_R3[4] DEC_Y_R3[5] DEC_Y_R3[6] 
+ DEC_Y_R3[7] DEC_Y_R4[0] DEC_Y_R4[1] DEC_Y_R4[2] DEC_Y_R4[3] DEC_Y_R4[4] 
+ DEC_Y_R4[5] DEC_Y_R4[6] DEC_Y_R4[7] S1AHSF400W40_SB_IO_SIM
XIO_LR AWT2_L2 AWT2_L1 BIST2IO_L2 BIST2IO_L1 BL_LR_1[0] BL_LR_1[1] BL_LR_1[2] 
+ BL_LR_1[3] BL_LR_1[4] BL_LR_1[5] BL_LR_1[6] BL_LR_1[7] BL_LR_1[8] BL_LR_1[9] 
+ BL_LR_1[10] BL_LR_1[11] BL_LR_1[12] BL_LR_1[13] BL_LR_1[14] BL_LR_1[15] 
+ BLB_LR_1[0] BLB_LR_1[1] BLB_LR_1[2] BLB_LR_1[3] BLB_LR_1[4] BLB_LR_1[5] 
+ BLB_LR_1[6] BLB_LR_1[7] BLB_LR_1[8] BLB_LR_1[9] BLB_LR_1[10] BLB_LR_1[11] 
+ BLB_LR_1[12] BLB_LR_1[13] BLB_LR_1[14] BLB_LR_1[15] BLEQ_L2 BLEQ_L1 BWEB_LR 
+ BWEBM_LR CKD_L2 CKD_L1 D_LR DM_LR PD_BUF_L2 PD_BUF_L1 Q_LR RE_L2 RE_L1 
+ SAE_L2 SAE_L1 VDDHD VDDI VSSI WE_L2 WE_L1 YL_L2[0] YL_L2[1] YL_L1[0] 
+ YL_L1[1] DEC_Y_L2[0] DEC_Y_L2[1] DEC_Y_L2[2] DEC_Y_L2[3] DEC_Y_L2[4] 
+ DEC_Y_L2[5] DEC_Y_L2[6] DEC_Y_L2[7] DEC_Y_L1[0] DEC_Y_L1[1] DEC_Y_L1[2] 
+ DEC_Y_L1[3] DEC_Y_L1[4] DEC_Y_L1[5] DEC_Y_L1[6] DEC_Y_L1[7] S1AHSF400W40_SB_IO_SIM
XIO_LL AWT2_L4 AWT2_L3 BIST2IO_L4 BIST2IO_L3 BL_LL_1[0] BL_LL_1[1] BL_LL_1[2] 
+ BL_LL_1[3] BL_LL_1[4] BL_LL_1[5] BL_LL_1[6] BL_LL_1[7] BL_LL_1[8] BL_LL_1[9] 
+ BL_LL_1[10] BL_LL_1[11] BL_LL_1[12] BL_LL_1[13] BL_LL_1[14] BL_LL_1[15] 
+ BLB_LL_1[0] BLB_LL_1[1] BLB_LL_1[2] BLB_LL_1[3] BLB_LL_1[4] BLB_LL_1[5] 
+ BLB_LL_1[6] BLB_LL_1[7] BLB_LL_1[8] BLB_LL_1[9] BLB_LL_1[10] BLB_LL_1[11] 
+ BLB_LL_1[12] BLB_LL_1[13] BLB_LL_1[14] BLB_LL_1[15] BLEQ_L4 BLEQ_L3 BWEB_LL 
+ BWEBM_LL CKD_L4 CKD_L3 D_LL DM_LL PD_BUF_L4 PD_BUF_L3 Q_LL RE_L4 RE_L3 
+ SAE_L4 SAE_L3 VDDHD VDDI VSSI WE_L4 WE_L3 YL_L4[0] YL_L4[1] YL_L3[0] 
+ YL_L3[1] DEC_Y_L4[0] DEC_Y_L4[1] DEC_Y_L4[2] DEC_Y_L4[3] DEC_Y_L4[4] 
+ DEC_Y_L4[5] DEC_Y_L4[6] DEC_Y_L4[7] DEC_Y_L3[0] DEC_Y_L3[1] DEC_Y_L3[2] 
+ DEC_Y_L3[3] DEC_Y_L3[4] DEC_Y_L3[5] DEC_Y_L3[6] DEC_Y_L3[7] S1AHSF400W40_SB_IO_SIM
XIO_RL AWT2_L1 AWT2_R2 BIST2IO_L1 BIST2IO_R2 NET0537[0] NET0537[1] NET0537[2] 
+ NET0537[3] NET0537[4] NET0537[5] NET0537[6] NET0537[7] NET0537[8] NET0537[9] 
+ NET0537[10] NET0537[11] NET0537[12] NET0537[13] NET0537[14] NET0537[15] 
+ NET0538[0] NET0538[1] NET0538[2] NET0538[3] NET0538[4] NET0538[5] NET0538[6] 
+ NET0538[7] NET0538[8] NET0538[9] NET0538[10] NET0538[11] NET0538[12] 
+ NET0538[13] NET0538[14] NET0538[15] BLEQ_L1 BLEQ_R2 NET0428 NET0360 CKD_L1 
+ CKD_R2 NET0534 NET0535 PD_BUF_L1 PD_BUF_R2 NET0361 RE_L1 RE_R2 SAE_L1 SAE_R2 
+ VDDHD VDDI VSSI WE_L1 WE_R2 YL_L1[0] YL_L1[1] YL_R2[0] YL_R2[1] DEC_Y_L1[0] 
+ DEC_Y_L1[1] DEC_Y_L1[2] DEC_Y_L1[3] DEC_Y_L1[4] DEC_Y_L1[5] DEC_Y_L1[6] 
+ DEC_Y_L1[7] DEC_Y_R2[0] DEC_Y_R2[1] DEC_Y_R2[2] DEC_Y_R2[3] DEC_Y_R2[4] 
+ DEC_Y_R2[5] DEC_Y_R2[6] DEC_Y_R2[7] S1AHSF400W40_SB_IO_SIM
XCNT AWT AWT2_L1 BIST BIST2IO_L1 BLEQ_L1 WL_TK CEB CEBM CKD_L1 CLK DEC_X0_1[0] 
+ DEC_X0_1[1] DEC_X0_1[2] DEC_X0_1[3] DEC_X0_1[4] DEC_X0_1[5] DEC_X0_1[6] 
+ DEC_X0_1[7] DEC_X1_1[0] DEC_X1_1[1] DEC_X1_1[2] DEC_X1_1[3] DEC_X1_1[4] 
+ DEC_X1_1[5] DEC_X1_1[6] DEC_X1_1[7] DEC_X2_1[0] DEC_X2_1[1] DEC_X2_1[2] 
+ DEC_X2_1[3] DEC_X2_1[4] DEC_X2_1[5] DEC_X2_1[6] DEC_X2_1[7] DEC_Y_L1[0] 
+ DEC_Y_L1[1] DEC_Y_L1[2] DEC_Y_L1[3] DEC_Y_L1[4] DEC_Y_L1[5] DEC_Y_L1[6] 
+ DEC_Y_L1[7] PD PD_BUF_L1 PTSEL RE_L1 RTSEL[0] RTSEL[1] SAE_L1 TK TM TRKBL 
+ VDDHD VDDI NET463 NET575 VSSI WE_L1 WEB WEBM WTSEL[0] WTSEL[1] WTSEL[2] X[0] 
+ X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] Y[0] Y[1] Y[2] Y[3] YL_L1[0] YL_L1[1] YM[0] YM[1] YM[2] 
+ YM[3] S1AHSF400W40_SB_CNT_SIM
XTKWL_LD VDDI TK_R2 TK_R3 VSSI WL_DUM_R2 WL_DUM_R3 WL_TK_R2 WL_TK_R3 
+ S1AHSF400W40_TKWL_LD_SIM
XTKWL_L VDDI TK TK_R2 VSSI WL_DUM_LT WL_DUM_R2 WL_TK WL_TK_R2 S1AHSF400W40_TKWL_SIM
XTKWL_R VDDI TK_R3 NET513 VSSI WL_DUM_R3 NET548 WL_TK_R3 WL_TK_LD S1AHSF400W40_TKWL_SIM
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_LCNT_M16_S64_U
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_LCNT_M16_S64_U BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] 
+ DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] 
+ DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] 
+ DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPYB_DN WLPYB_UP 
+ WLPY_DN WLPY_UP WLP_SAE WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO BLEQ_DN:B BLEQ_UP:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B DEC_Y_DN[0]:B DEC_Y_DN[1]:B DEC_Y_DN[2]:B DEC_Y_DN[3]:B 
*.PININFO DEC_Y_DN[4]:B DEC_Y_DN[5]:B DEC_Y_DN[6]:B DEC_Y_DN[7]:B 
*.PININFO DEC_Y_UP[0]:B DEC_Y_UP[1]:B DEC_Y_UP[2]:B DEC_Y_UP[3]:B 
*.PININFO DEC_Y_UP[4]:B DEC_Y_UP[5]:B DEC_Y_UP[6]:B DEC_Y_UP[7]:B PD_BUF:B 
*.PININFO RE:B RW_RE:B SAEB:B VDDHD:B VDDI:B VSSI:B WE:B WLPYB_DN:B WLPYB_UP:B 
*.PININFO WLPY_DN:B WLPY_UP:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B YL_LIO[0]:B 
*.PININFO YL_LIO[1]:B
XLCNT BLEQ_DN BLEQ_UP NET049[0] NET049[1] NET049[2] NET049[3] NET049[4] 
+ NET049[5] NET049[6] NET049[7] NET048[0] NET048[1] NET048[2] NET048[3] 
+ NET048[4] NET048[5] NET048[6] NET048[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[6] DEC_X3[7] NET045[0] NET045[1] NET045[2] NET045[3] 
+ NET045[4] NET045[5] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF NET46 RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN WLPY_1[1] WLPY_1[2] 
+ WLPY_1[3] WLPY_UP WLPY_2[1] WLPY_2[2] WLPY_2[3] WLP_SAE NET010 YL[0] 
+ YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL_F_M16
XI3 VDDHD VDDI VSSI WLPY_UP WLPYB_UP S1AHSF400W40_XDRV_STRAP
XXDRV_STRP VDDHD VDDI VSSI WLPY_DN WLPYB_DN S1AHSF400W40_XDRV_STRAP
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_LCNT_M8_S64_U
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_LCNT_M8_S64_U BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] 
+ DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] 
+ DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] 
+ DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPYB_DN WLPYB_UP 
+ WLPY_DN WLPY_UP WLP_SAE WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO BLEQ_DN:B BLEQ_UP:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B DEC_Y_DN[0]:B DEC_Y_DN[1]:B DEC_Y_DN[2]:B DEC_Y_DN[3]:B 
*.PININFO DEC_Y_DN[4]:B DEC_Y_DN[5]:B DEC_Y_DN[6]:B DEC_Y_DN[7]:B 
*.PININFO DEC_Y_UP[0]:B DEC_Y_UP[1]:B DEC_Y_UP[2]:B DEC_Y_UP[3]:B 
*.PININFO DEC_Y_UP[4]:B DEC_Y_UP[5]:B DEC_Y_UP[6]:B DEC_Y_UP[7]:B PD_BUF:B 
*.PININFO RE:B RW_RE:B SAEB:B VDDHD:B VDDI:B VSSI:B WE:B WLPYB_DN:B WLPYB_UP:B 
*.PININFO WLPY_DN:B WLPY_UP:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B YL_LIO[0]:B 
*.PININFO YL_LIO[1]:B
XLCNT BLEQ_DN BLEQ_UP NET049[0] NET049[1] NET049[2] NET049[3] NET049[4] 
+ NET049[5] NET049[6] NET049[7] NET048[0] NET048[1] NET048[2] NET048[3] 
+ NET048[4] NET048[5] NET048[6] NET048[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[6] DEC_X3[7] NET046[0] NET046[1] NET046[2] NET046[3] 
+ NET046[4] NET046[5] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF NET46 RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN WLPY_1[1] WLPY_1[2] 
+ WLPY_1[3] WLPY_UP WLPY_2[1] WLPY_2[2] WLPY_2[3] WLP_SAE NET045 YL[0] 
+ YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL_F_M8
XI3 VDDHD VDDI VSSI WLPY_UP WLPYB_UP S1AHSF400W40_XDRV_STRAP
XXDRV_STRP VDDHD VDDI VSSI WLPY_DN WLPYB_DN S1AHSF400W40_XDRV_STRAP
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_LCNT_M4_S64_U
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_LCNT_M4_S64_U BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] 
+ DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] 
+ DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] 
+ DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPYB_DN WLPYB_UP 
+ WLPY_DN WLPY_UP WLP_SAE WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO BLEQ_DN:B BLEQ_UP:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B DEC_Y_DN[0]:B DEC_Y_DN[1]:B DEC_Y_DN[2]:B DEC_Y_DN[3]:B 
*.PININFO DEC_Y_DN[4]:B DEC_Y_DN[5]:B DEC_Y_DN[6]:B DEC_Y_DN[7]:B 
*.PININFO DEC_Y_UP[0]:B DEC_Y_UP[1]:B DEC_Y_UP[2]:B DEC_Y_UP[3]:B 
*.PININFO DEC_Y_UP[4]:B DEC_Y_UP[5]:B DEC_Y_UP[6]:B DEC_Y_UP[7]:B PD_BUF:B 
*.PININFO RE:B RW_RE:B SAEB:B VDDHD:B VDDI:B VSSI:B WE:B WLPYB_DN:B WLPYB_UP:B 
*.PININFO WLPY_DN:B WLPY_UP:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B YL_LIO[0]:B 
*.PININFO YL_LIO[1]:B
XLCNT BLEQ_DN BLEQ_UP NET049[0] NET049[1] NET049[2] NET049[3] NET049[4] 
+ NET049[5] NET049[6] NET049[7] NET048[0] NET048[1] NET048[2] NET048[3] 
+ NET048[4] NET048[5] NET048[6] NET048[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[6] DEC_X3[7] NET046[0] NET046[1] NET046[2] NET046[3] 
+ NET046[4] NET046[5] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF NET46 RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN WLPY_1[1] WLPY_1[2] 
+ WLPY_1[3] WLPY_UP WLPY_2[1] WLPY_2[2] WLPY_2[3] WLP_SAE NET045 YL[0] 
+ YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL_F_M4
XI3 VDDHD VDDI VSSI WLPY_UP WLPYB_UP S1AHSF400W40_XDRV_STRAP
XXDRV_STRP VDDHD VDDI VSSI WLPY_DN WLPYB_DN S1AHSF400W40_XDRV_STRAP
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_LCNT_M8_S256_U
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_LCNT_M8_S256_U BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] 
+ DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] 
+ DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] 
+ DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPYB_DN WLPYB_UP 
+ WLPY_DN WLPY_UP WLP_SAE WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO BLEQ_DN:B BLEQ_UP:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B DEC_Y_DN[0]:B DEC_Y_DN[1]:B DEC_Y_DN[2]:B DEC_Y_DN[3]:B 
*.PININFO DEC_Y_DN[4]:B DEC_Y_DN[5]:B DEC_Y_DN[6]:B DEC_Y_DN[7]:B 
*.PININFO DEC_Y_UP[0]:B DEC_Y_UP[1]:B DEC_Y_UP[2]:B DEC_Y_UP[3]:B 
*.PININFO DEC_Y_UP[4]:B DEC_Y_UP[5]:B DEC_Y_UP[6]:B DEC_Y_UP[7]:B PD_BUF:B 
*.PININFO RE:B RW_RE:B SAEB:B VDDHD:B VDDI:B VSSI:B WE:B WLPYB_DN:B WLPYB_UP:B 
*.PININFO WLPY_DN:B WLPY_UP:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B YL_LIO[0]:B 
*.PININFO YL_LIO[1]:B
XLCNT BLEQ_DN BLEQ_UP NET045[0] NET045[1] NET045[2] NET045[3] NET045[4] 
+ NET045[5] NET045[6] NET045[7] NET046[0] NET046[1] NET046[2] NET046[3] 
+ NET046[4] NET046[5] NET046[6] NET046[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[6] DEC_X3[7] NET049[0] NET049[1] NET049[2] NET049[3] 
+ NET049[4] NET049[5] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF NET46 RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN WLPY_1[1] WLPY_1[2] 
+ WLPY_1[3] WLPY_2[0] WLPY_2[1] WLPY_2[2] WLPY_UP WLP_SAE NET010 YL[0] 
+ YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL_S_M8
XI3 VDDHD VDDI VSSI WLPY_UP WLPYB_UP S1AHSF400W40_XDRV_STRAP
XXDRV_STRP VDDHD VDDI VSSI WLPY_DN WLPYB_DN S1AHSF400W40_XDRV_STRAP
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_LCNT_M16_S256_U
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_LCNT_M16_S256_U BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] 
+ DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] 
+ DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] 
+ DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPYB_DN WLPYB_UP 
+ WLPY_DN WLPY_UP WLP_SAE WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO BLEQ_DN:B BLEQ_UP:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B DEC_Y_DN[0]:B DEC_Y_DN[1]:B DEC_Y_DN[2]:B DEC_Y_DN[3]:B 
*.PININFO DEC_Y_DN[4]:B DEC_Y_DN[5]:B DEC_Y_DN[6]:B DEC_Y_DN[7]:B 
*.PININFO DEC_Y_UP[0]:B DEC_Y_UP[1]:B DEC_Y_UP[2]:B DEC_Y_UP[3]:B 
*.PININFO DEC_Y_UP[4]:B DEC_Y_UP[5]:B DEC_Y_UP[6]:B DEC_Y_UP[7]:B PD_BUF:B 
*.PININFO RE:B RW_RE:B SAEB:B VDDHD:B VDDI:B VSSI:B WE:B WLPYB_DN:B WLPYB_UP:B 
*.PININFO WLPY_DN:B WLPY_UP:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B YL_LIO[0]:B 
*.PININFO YL_LIO[1]:B
XLCNT BLEQ_DN BLEQ_UP NET049[0] NET049[1] NET049[2] NET049[3] NET049[4] 
+ NET049[5] NET049[6] NET049[7] NET045[0] NET045[1] NET045[2] NET045[3] 
+ NET045[4] NET045[5] NET045[6] NET045[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[6] DEC_X3[7] NET048[0] NET048[1] NET048[2] NET048[3] 
+ NET048[4] NET048[5] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF NET46 RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN WLPY_1[1] WLPY_1[2] 
+ WLPY_1[3] WLPY_2[0] WLPY_2[1] WLPY_2[2] WLPY_UP WLP_SAE NET010 YL[0] 
+ YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL_S_M16
XI3 VDDHD VDDI VSSI WLPY_UP WLPYB_UP S1AHSF400W40_XDRV_STRAP
XXDRV_STRP VDDHD VDDI VSSI WLPY_DN WLPYB_DN S1AHSF400W40_XDRV_STRAP
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_LCNT_M4_S256_U
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_LCNT_M4_S256_U BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] 
+ DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] 
+ DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] 
+ DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] 
+ DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] 
+ DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] 
+ DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPYB_DN WLPYB_UP 
+ WLPY_DN WLPY_UP WLP_SAE WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO BLEQ_DN:B BLEQ_UP:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B DEC_Y_DN[0]:B DEC_Y_DN[1]:B DEC_Y_DN[2]:B DEC_Y_DN[3]:B 
*.PININFO DEC_Y_DN[4]:B DEC_Y_DN[5]:B DEC_Y_DN[6]:B DEC_Y_DN[7]:B 
*.PININFO DEC_Y_UP[0]:B DEC_Y_UP[1]:B DEC_Y_UP[2]:B DEC_Y_UP[3]:B 
*.PININFO DEC_Y_UP[4]:B DEC_Y_UP[5]:B DEC_Y_UP[6]:B DEC_Y_UP[7]:B PD_BUF:B 
*.PININFO RE:B RW_RE:B SAEB:B VDDHD:B VDDI:B VSSI:B WE:B WLPYB_DN:B WLPYB_UP:B 
*.PININFO WLPY_DN:B WLPY_UP:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B YL_LIO[0]:B 
*.PININFO YL_LIO[1]:B
XI3 VDDHD VDDI VSSI WLPY_UP WLPYB_UP S1AHSF400W40_XDRV_STRAP
XXDRV_STRP VDDHD VDDI VSSI WLPY_DN WLPYB_DN S1AHSF400W40_XDRV_STRAP
XLCNT BLEQ_DN BLEQ_UP NET060[0] NET060[1] NET060[2] NET060[3] NET060[4] 
+ NET060[5] NET060[6] NET060[7] NET061[0] NET061[1] NET061[2] NET061[3] 
+ NET061[4] NET061[5] NET061[6] NET061[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[6] DEC_X3[7] NET059[0] NET059[1] NET059[2] NET059[3] 
+ NET059[4] NET059[5] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF NET46 RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN WLPY_1[1] WLPY_1[2] 
+ WLPY_1[3] WLPY_2[0] WLPY_2[1] WLPY_2[2] WLPY_UP WLP_SAE NET057 YL[0] 
+ YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL_S_M4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_LCNT_U_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_LCNT_U_SIM BLEQ_DN_LT BLEQ_DN_RT BLEQ_UP_LT BLEQ_UP_RT CVDDHD CVDDI 
+ DEC_X0_BT[0] DEC_X0_BT[1] DEC_X0_BT[2] DEC_X0_BT[3] DEC_X0_BT[4] 
+ DEC_X0_BT[5] DEC_X0_BT[6] DEC_X0_BT[7] DEC_X0_TP[0] DEC_X0_TP[1] 
+ DEC_X0_TP[2] DEC_X0_TP[3] DEC_X0_TP[4] DEC_X0_TP[5] DEC_X0_TP[6] 
+ DEC_X0_TP[7] DEC_X1_BT[0] DEC_X1_BT[1] DEC_X1_BT[2] DEC_X1_BT[3] 
+ DEC_X1_BT[4] DEC_X1_BT[5] DEC_X1_BT[6] DEC_X1_BT[7] DEC_X1_TP[0] 
+ DEC_X1_TP[1] DEC_X1_TP[2] DEC_X1_TP[3] DEC_X1_TP[4] DEC_X1_TP[5] 
+ DEC_X1_TP[6] DEC_X1_TP[7] DEC_X2_BT[0] DEC_X2_BT[1] DEC_X2_BT[2] 
+ DEC_X2_BT[3] DEC_X2_TP[0] DEC_X2_TP[1] DEC_X2_TP[2] DEC_X2_TP[3] 
+ DEC_X3_BT[0] DEC_X3_BT[1] DEC_X3_BT[2] DEC_X3_BT[3] DEC_X3_BT[4] 
+ DEC_X3_BT[5] DEC_X3_BT[6] DEC_X3_BT[7] DEC_X3_TP[0] DEC_X3_TP[1] 
+ DEC_X3_TP[2] DEC_X3_TP[3] DEC_X3_TP[4] DEC_X3_TP[5] DEC_X3_TP[6] 
+ DEC_X3_TP[7] DEC_Y_BT[0] DEC_Y_BT[1] DEC_Y_BT[2] DEC_Y_BT[3] DEC_Y_BT[4] 
+ DEC_Y_BT[5] DEC_Y_BT[6] DEC_Y_BT[7] DEC_Y_DN_LT[0] DEC_Y_DN_LT[1] 
+ DEC_Y_DN_LT[2] DEC_Y_DN_LT[3] DEC_Y_DN_LT[4] DEC_Y_DN_LT[5] DEC_Y_DN_LT[6] 
+ DEC_Y_DN_LT[7] DEC_Y_DN_RT[0] DEC_Y_DN_RT[1] DEC_Y_DN_RT[2] DEC_Y_DN_RT[3] 
+ DEC_Y_DN_RT[4] DEC_Y_DN_RT[5] DEC_Y_DN_RT[6] DEC_Y_DN_RT[7] DEC_Y_TP[0] 
+ DEC_Y_TP[1] DEC_Y_TP[2] DEC_Y_TP[3] DEC_Y_TP[4] DEC_Y_TP[5] DEC_Y_TP[6] 
+ DEC_Y_TP[7] DEC_Y_UP_LT[0] DEC_Y_UP_LT[1] DEC_Y_UP_LT[2] DEC_Y_UP_LT[3] 
+ DEC_Y_UP_LT[4] DEC_Y_UP_LT[5] DEC_Y_UP_LT[6] DEC_Y_UP_LT[7] DEC_Y_UP_RT[0] 
+ DEC_Y_UP_RT[1] DEC_Y_UP_RT[2] DEC_Y_UP_RT[3] DEC_Y_UP_RT[4] DEC_Y_UP_RT[5] 
+ DEC_Y_UP_RT[6] DEC_Y_UP_RT[7] PD_BUF_BT PD_BUF_TP PD_CVDDBUF_BT 
+ PD_CVDDBUF_TP RE_LT RE_RT RW_RE_BT RW_RE_TP SAEB_LT SAEB_RT VDDHD VDDI VSSI 
+ WE_LT WE_RT WLPYB_DN_BT WLPYB_UP_TP WLPY_DN_BT WLPY_UP_TP WLP_SAE_BT 
+ WLP_SAE_TK_BT WLP_SAE_TK_TP WLP_SAE_TP YL_BT[0] YL_LIO_LT[0] YL_LIO_LT[1] 
+ YL_LIO_RT[0] YL_LIO_RT[1] YL_TP[0]
*.PININFO DEC_X0_BT[0]:I DEC_X0_BT[1]:I DEC_X0_BT[2]:I DEC_X0_BT[3]:I 
*.PININFO DEC_X0_BT[4]:I DEC_X0_BT[5]:I DEC_X0_BT[6]:I DEC_X0_BT[7]:I 
*.PININFO DEC_X1_BT[0]:I DEC_X1_BT[1]:I DEC_X1_BT[2]:I DEC_X1_BT[3]:I 
*.PININFO DEC_X1_BT[4]:I DEC_X1_BT[5]:I DEC_X1_BT[6]:I DEC_X1_BT[7]:I 
*.PININFO PD_BUF_BT:I PD_CVDDBUF_BT:I RW_RE_TP:I DEC_X0_TP[0]:O DEC_X0_TP[1]:O 
*.PININFO DEC_X0_TP[2]:O DEC_X0_TP[3]:O DEC_X0_TP[4]:O DEC_X0_TP[5]:O 
*.PININFO DEC_X0_TP[6]:O DEC_X0_TP[7]:O DEC_X1_TP[0]:O DEC_X1_TP[1]:O 
*.PININFO DEC_X1_TP[2]:O DEC_X1_TP[3]:O DEC_X1_TP[4]:O DEC_X1_TP[5]:O 
*.PININFO DEC_X1_TP[6]:O DEC_X1_TP[7]:O PD_BUF_TP:O PD_CVDDBUF_TP:O 
*.PININFO BLEQ_DN_LT:B BLEQ_DN_RT:B BLEQ_UP_LT:B BLEQ_UP_RT:B CVDDHD:B CVDDI:B 
*.PININFO DEC_X2_BT[0]:B DEC_X2_BT[1]:B DEC_X2_BT[2]:B DEC_X2_BT[3]:B 
*.PININFO DEC_X2_TP[0]:B DEC_X2_TP[1]:B DEC_X2_TP[2]:B DEC_X2_TP[3]:B 
*.PININFO DEC_X3_BT[0]:B DEC_X3_BT[1]:B DEC_X3_BT[2]:B DEC_X3_BT[3]:B 
*.PININFO DEC_X3_BT[4]:B DEC_X3_BT[5]:B DEC_X3_BT[6]:B DEC_X3_BT[7]:B 
*.PININFO DEC_X3_TP[0]:B DEC_X3_TP[1]:B DEC_X3_TP[2]:B DEC_X3_TP[3]:B 
*.PININFO DEC_X3_TP[4]:B DEC_X3_TP[5]:B DEC_X3_TP[6]:B DEC_X3_TP[7]:B 
*.PININFO DEC_Y_BT[0]:B DEC_Y_BT[1]:B DEC_Y_BT[2]:B DEC_Y_BT[3]:B 
*.PININFO DEC_Y_BT[4]:B DEC_Y_BT[5]:B DEC_Y_BT[6]:B DEC_Y_BT[7]:B 
*.PININFO DEC_Y_DN_LT[0]:B DEC_Y_DN_LT[1]:B DEC_Y_DN_LT[2]:B DEC_Y_DN_LT[3]:B 
*.PININFO DEC_Y_DN_LT[4]:B DEC_Y_DN_LT[5]:B DEC_Y_DN_LT[6]:B DEC_Y_DN_LT[7]:B 
*.PININFO DEC_Y_DN_RT[0]:B DEC_Y_DN_RT[1]:B DEC_Y_DN_RT[2]:B DEC_Y_DN_RT[3]:B 
*.PININFO DEC_Y_DN_RT[4]:B DEC_Y_DN_RT[5]:B DEC_Y_DN_RT[6]:B DEC_Y_DN_RT[7]:B 
*.PININFO DEC_Y_TP[0]:B DEC_Y_TP[1]:B DEC_Y_TP[2]:B DEC_Y_TP[3]:B 
*.PININFO DEC_Y_TP[4]:B DEC_Y_TP[5]:B DEC_Y_TP[6]:B DEC_Y_TP[7]:B 
*.PININFO DEC_Y_UP_LT[0]:B DEC_Y_UP_LT[1]:B DEC_Y_UP_LT[2]:B DEC_Y_UP_LT[3]:B 
*.PININFO DEC_Y_UP_LT[4]:B DEC_Y_UP_LT[5]:B DEC_Y_UP_LT[6]:B DEC_Y_UP_LT[7]:B 
*.PININFO DEC_Y_UP_RT[0]:B DEC_Y_UP_RT[1]:B DEC_Y_UP_RT[2]:B DEC_Y_UP_RT[3]:B 
*.PININFO DEC_Y_UP_RT[4]:B DEC_Y_UP_RT[5]:B DEC_Y_UP_RT[6]:B DEC_Y_UP_RT[7]:B 
*.PININFO RE_LT:B RE_RT:B RW_RE_BT:B SAEB_LT:B SAEB_RT:B VDDHD:B VDDI:B VSSI:B 
*.PININFO WE_LT:B WE_RT:B WLPYB_DN_BT:B WLPYB_UP_TP:B WLPY_DN_BT:B 
*.PININFO WLPY_UP_TP:B WLP_SAE_BT:B WLP_SAE_TK_BT:B WLP_SAE_TK_TP:B 
*.PININFO WLP_SAE_TP:B YL_BT[0]:B YL_LIO_LT[0]:B YL_LIO_LT[1]:B YL_LIO_RT[0]:B 
*.PININFO YL_LIO_RT[1]:B YL_TP[0]:B
XI26 NET080 NET079 NET078[0] NET078[1] NET078[2] NET078[3] NET078[4] NET078[5] 
+ NET078[6] NET078[7] NET077[0] NET077[1] NET077[2] NET077[3] NET077[4] 
+ NET077[5] NET077[6] NET077[7] NET076[0] NET076[1] NET076[2] NET076[3] 
+ NET012[0] NET012[1] NET012[2] NET012[3] NET012[4] NET012[5] NET012[6] 
+ NET012[7] NET074[0] NET074[1] NET074[2] NET074[3] NET074[4] NET074[5] 
+ NET074[6] NET074[7] NET073[0] NET073[1] NET073[2] NET073[3] NET073[4] 
+ NET073[5] NET073[6] NET073[7] NET05[0] NET05[1] NET05[2] NET05[3] NET05[4] 
+ NET05[5] NET05[6] NET05[7] NET010 NET09 NET015 NET018 NET04 NET03 NET016 
+ NET014 NET083 NET082 NET08 NET06 NET017 NET081 NET07 NET011[0] NET011[1] 
+ S1AHSF400W40_BK_LCNT_M16_S64_U
XI25 NET0105 NET0104 NET0103[0] NET0103[1] NET0103[2] NET0103[3] NET0103[4] 
+ NET0103[5] NET0103[6] NET0103[7] NET0102[0] NET0102[1] NET0102[2] NET0102[3] 
+ NET0102[4] NET0102[5] NET0102[6] NET0102[7] NET0101[0] NET0101[1] NET0101[2] 
+ NET0101[3] NET0100[0] NET0100[1] NET0100[2] NET0100[3] NET0100[4] NET0100[5] 
+ NET0100[6] NET0100[7] NET099[0] NET099[1] NET099[2] NET099[3] NET099[4] 
+ NET099[5] NET099[6] NET099[7] NET098[0] NET098[1] NET098[2] NET098[3] 
+ NET098[4] NET098[5] NET098[6] NET098[7] NET097[0] NET097[1] NET097[2] 
+ NET097[3] NET097[4] NET097[5] NET097[6] NET097[7] NET096 NET095 NET094 
+ NET093 NET092 NET091 NET090 NET089 NET0108 NET0107 NET088 NET087 NET086 
+ NET0106 NET085 NET084[0] NET084[1] S1AHSF400W40_BK_LCNT_M8_S64_U
XI27 NET0130 NET0129 NET0128[0] NET0128[1] NET0128[2] NET0128[3] NET0128[4] 
+ NET0128[5] NET0128[6] NET0128[7] NET0127[0] NET0127[1] NET0127[2] NET0127[3] 
+ NET0127[4] NET0127[5] NET0127[6] NET0127[7] NET0126[0] NET0126[1] NET0126[2] 
+ NET0126[3] NET0125[0] NET0125[1] NET0125[2] NET0125[3] NET0125[4] NET0125[5] 
+ NET0125[6] NET0125[7] NET0124[0] NET0124[1] NET0124[2] NET0124[3] NET0124[4] 
+ NET0124[5] NET0124[6] NET0124[7] NET0123[0] NET0123[1] NET0123[2] NET0123[3] 
+ NET0123[4] NET0123[5] NET0123[6] NET0123[7] NET0122[0] NET0122[1] NET0122[2] 
+ NET0122[3] NET0122[4] NET0122[5] NET0122[6] NET0122[7] NET0121 NET0120 
+ NET0119 NET0118 NET0117 NET0116 NET0115 NET0114 NET0133 NET0132 NET0113 
+ NET0112 NET0111 NET0131 NET0110 NET0109[0] NET0109[1] S1AHSF400W40_BK_LCNT_M4_S64_U
XI23 NET069 NET068 NET067[0] NET067[1] NET067[2] NET067[3] NET067[4] NET067[5] 
+ NET067[6] NET067[7] NET066[0] NET066[1] NET066[2] NET066[3] NET066[4] 
+ NET066[5] NET066[6] NET066[7] NET065[0] NET065[1] NET065[2] NET065[3] 
+ NET064[0] NET064[1] NET064[2] NET064[3] NET064[4] NET064[5] NET064[6] 
+ NET064[7] NET063[0] NET063[1] NET063[2] NET063[3] NET063[4] NET063[5] 
+ NET063[6] NET063[7] NET062[0] NET062[1] NET062[2] NET062[3] NET062[4] 
+ NET062[5] NET062[6] NET062[7] NET061[0] NET061[1] NET061[2] NET061[3] 
+ NET061[4] NET061[5] NET061[6] NET061[7] NET060 NET059 NET058 NET057 NET056 
+ NET055 NET054 NET053 NET071 NET070 NET052 NET051 NET050 NET013 NET01 
+ NET02[0] NET02[1] S1AHSF400W40_BK_LCNT_M8_S256_U
XI24 NET0180 NET0179 NET0178[0] NET0178[1] NET0178[2] NET0178[3] NET0178[4] 
+ NET0178[5] NET0178[6] NET0178[7] NET0177[0] NET0177[1] NET0177[2] NET0177[3] 
+ NET0177[4] NET0177[5] NET0177[6] NET0177[7] NET0176[0] NET0176[1] NET0176[2] 
+ NET0176[3] NET0175[0] NET0175[1] NET0175[2] NET0175[3] NET0175[4] NET0175[5] 
+ NET0175[6] NET0175[7] NET0174[0] NET0174[1] NET0174[2] NET0174[3] NET0174[4] 
+ NET0174[5] NET0174[6] NET0174[7] NET0173[0] NET0173[1] NET0173[2] NET0173[3] 
+ NET0173[4] NET0173[5] NET0173[6] NET0173[7] NET0172[0] NET0172[1] NET0172[2] 
+ NET0172[3] NET0172[4] NET0172[5] NET0172[6] NET0172[7] NET0171 NET0170 
+ NET0169 NET0168 NET0167 NET0166 NET0165 NET0164 NET0183 NET0182 NET0163 
+ NET0162 NET0161 NET0181 NET0160 NET0159[0] NET0159[1] S1AHSF400W40_BK_LCNT_M16_S256_U
XI22 NET68 NET67 NET66[0] NET66[1] NET66[2] NET66[3] NET66[4] NET66[5] 
+ NET66[6] NET66[7] NET65[0] NET65[1] NET65[2] NET65[3] NET65[4] NET65[5] 
+ NET65[6] NET65[7] NET64[0] NET64[1] NET64[2] NET64[3] NET63[0] NET63[1] 
+ NET63[2] NET63[3] NET63[4] NET63[5] NET63[6] NET63[7] NET62[0] NET62[1] 
+ NET62[2] NET62[3] NET62[4] NET62[5] NET62[6] NET62[7] NET61[0] NET61[1] 
+ NET61[2] NET61[3] NET61[4] NET61[5] NET61[6] NET61[7] NET60[0] NET60[1] 
+ NET60[2] NET60[3] NET60[4] NET60[5] NET60[6] NET60[7] NET59 NET57 NET56 
+ NET55 NET54 NET53 NET52 NET51 NET049 NET048 NET047 NET046 NET48 NET075 
+ NET072 NET46[0] NET46[1] S1AHSF400W40_BK_LCNT_M4_S256_U
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    ARR_LIO2_SEG6_S64
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ARR_LIO2_SEG6_S64 CVDDI GBL GBLB GW GWB VDDHD VDDI VSSI
*.PININFO CVDDI:B GBL:B GBLB:B GW:B GWB:B VDDHD:B VDDI:B VSSI:B
XI39 NET053[0] NET053[1] NET053[2] NET053[3] NET052[0] NET052[1] NET052[2] 
+ NET052[3] GBL GBLB GW GWB VDDI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI S1AHSF400W40_MCB_64X4_CHAR
XI34 BL_UP_1[0] BL_UP_1[1] BL_UP_1[2] BL_UP_1[3] BLB_UP_1[0] BLB_UP_1[1] 
+ BLB_UP_1[2] BLB_UP_1[3] GBL GBLB GW GWB VDDI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ S1AHSF400W40_MCB_64X4_CHAR
XI36 BL_DN_0[0] BL_DN_0[1] BL_DN_0[2] BL_DN_0[3] BLB_DN_0[0] BLB_DN_0[1] 
+ BLB_DN_0[2] BLB_DN_0[3] GBL GBLB GW GWB VDDI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ S1AHSF400W40_MCB_64X4_CHAR
XI35 BL_UP_0[0] BL_UP_0[1] BL_UP_0[2] BL_UP_0[3] BLB_UP_0[0] BLB_UP_0[1] 
+ BLB_UP_0[2] BLB_UP_0[3] GBL GBLB GW GWB VDDI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ S1AHSF400W40_MCB_64X4_CHAR
XI38 NET071[0] NET071[1] NET071[2] NET071[3] NET070[0] NET070[1] NET070[2] 
+ NET070[3] GBL GBLB GW GWB VDDI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI S1AHSF400W40_MCB_64X4_CHAR
XI33 BL_DN_1[0] BL_DN_1[1] BL_DN_1[2] BL_DN_1[3] BLB_DN_1[0] BLB_DN_1[1] 
+ BLB_DN_1[2] BLB_DN_1[3] GBL GBLB GW GWB VDDI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ S1AHSF400W40_MCB_64X4_CHAR
XLIO_M4 BLB_DN_1[0] BLB_DN_1[1] BLB_DN_1[2] BLB_DN_1[3] BLB_UP_1[0] 
+ BLB_UP_1[1] BLB_UP_1[2] BLB_UP_1[3] VDDI VDDI BL_DN_1[0] BL_DN_1[1] 
+ BL_DN_1[2] BL_DN_1[3] BL_UP_1[0] BL_UP_1[1] BL_UP_1[2] BL_UP_1[3] GBL GBLB 
+ GW GWB VSSI VDDI VDDHD VDDI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI S1AHSF400W40_LIO_M4
XI37 BLB_DN_0[0] BLB_DN_0[1] BLB_DN_0[2] BLB_DN_0[3] BLB_UP_0[0] BLB_UP_0[1] 
+ BLB_UP_0[2] BLB_UP_0[3] VDDI VDDI BL_DN_0[0] BL_DN_0[1] BL_DN_0[2] 
+ BL_DN_0[3] BL_UP_0[0] BL_UP_0[1] BL_UP_0[2] BL_UP_0[3] GBL GBLB GW GWB VSSI 
+ VDDI VDDHD VDDI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI S1AHSF400W40_LIO_M4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    ARR_LIO2_SEG6_S256
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ARR_LIO2_SEG6_S256 CVDDI GBL GBLB GW GWB VDDHD VDDI VSSI
*.PININFO CVDDI:B GBL:B GBLB:B GW:B GWB:B VDDHD:B VDDI:B VSSI:B
XI39 NET053[0] NET053[1] NET053[2] NET053[3] NET052[0] NET052[1] NET052[2] 
+ NET052[3] GBL GBLB GW GWB VDDI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI S1AHSF400W40_MCB_256X4_CHAR
XI34 BL_UP_1[0] BL_UP_1[1] BL_UP_1[2] BL_UP_1[3] BLB_UP_1[0] BLB_UP_1[1] 
+ BLB_UP_1[2] BLB_UP_1[3] GBL GBLB GW GWB VDDI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI S1AHSF400W40_MCB_256X4_CHAR
XI36 BL_DN_0[0] BL_DN_0[1] BL_DN_0[2] BL_DN_0[3] BLB_DN_0[0] BLB_DN_0[1] 
+ BLB_DN_0[2] BLB_DN_0[3] GBL GBLB GW GWB VDDI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI S1AHSF400W40_MCB_256X4_CHAR
XI35 BL_UP_0[0] BL_UP_0[1] BL_UP_0[2] BL_UP_0[3] BLB_UP_0[0] BLB_UP_0[1] 
+ BLB_UP_0[2] BLB_UP_0[3] GBL GBLB GW GWB VDDI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI S1AHSF400W40_MCB_256X4_CHAR
XI38 NET071[0] NET071[1] NET071[2] NET071[3] NET070[0] NET070[1] NET070[2] 
+ NET070[3] GBL GBLB GW GWB VDDI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI S1AHSF400W40_MCB_256X4_CHAR
XI33 BL_DN_1[0] BL_DN_1[1] BL_DN_1[2] BL_DN_1[3] BLB_DN_1[0] BLB_DN_1[1] 
+ BLB_DN_1[2] BLB_DN_1[3] GBL GBLB GW GWB VDDI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI S1AHSF400W40_MCB_256X4_CHAR
XLIO_M4 BLB_DN_1[0] BLB_DN_1[1] BLB_DN_1[2] BLB_DN_1[3] BLB_UP_1[0] 
+ BLB_UP_1[1] BLB_UP_1[2] BLB_UP_1[3] VDDI VDDI BL_DN_1[0] BL_DN_1[1] 
+ BL_DN_1[2] BL_DN_1[3] BL_UP_1[0] BL_UP_1[1] BL_UP_1[2] BL_UP_1[3] GBL GBLB 
+ GW GWB VSSI VDDI VDDHD VDDI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI S1AHSF400W40_LIO_M4
XI37 BLB_DN_0[0] BLB_DN_0[1] BLB_DN_0[2] BLB_DN_0[3] BLB_UP_0[0] BLB_UP_0[1] 
+ BLB_UP_0[2] BLB_UP_0[3] VDDI VDDI BL_DN_0[0] BL_DN_0[1] BL_DN_0[2] 
+ BL_DN_0[3] BL_UP_0[0] BL_UP_0[1] BL_UP_0[2] BL_UP_0[3] GBL GBLB GW GWB VSSI 
+ VDDI VDDHD VDDI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI S1AHSF400W40_LIO_M4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    ARR_SEG_LD_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ARR_SEG_LD_SIM CVDDI GBLB_BT GBLB_TP GBL_BT GBL_TP GWB_BT GWB_TP GW_BT 
+ GW_TP VDDHD VDDI VSSI
*.PININFO CVDDI:B GBLB_BT:B GBLB_TP:B GBL_BT:B GBL_TP:B GWB_BT:B GWB_TP:B 
*.PININFO GW_BT:B GW_TP:B VDDHD:B VDDI:B VSSI:B
XI34 NET016 NET017 NET015 NET014 NET013 NET020 NET019 NET018 
+ S1AHSF400W40_ARR_LIO2_SEG6_S64
XI33 NET17 NET16 NET15 NET14 NET13 NET20 NET19 NET18 S1AHSF400W40_ARR_LIO2_SEG6_S256
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_LCNT2_SEG6_S64
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_LCNT2_SEG6_S64 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] 
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] PD_BUF RW_RE VDDHD VDDI VSSI WLP_SAE WLP_SAE_TK YL[0]
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B DEC_X3[4]:B 
*.PININFO DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B DEC_Y[1]:B DEC_Y[2]:B 
*.PININFO DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B DEC_Y[7]:B PD_BUF:B 
*.PININFO RW_RE:B VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XI4 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] PD_BUF PD_CVDDBUF VDDHD VDDI VSSI NET39[0] NET39[1] 
+ NET39[2] NET39[3] NET39[4] NET39[5] NET39[6] NET39[7] NET39[8] NET39[9] 
+ NET39[10] NET39[11] NET39[12] NET39[13] NET39[14] NET39[15] NET39[16] 
+ NET39[17] NET39[18] NET39[19] NET39[20] NET39[21] NET39[22] NET39[23] 
+ NET39[24] NET39[25] NET39[26] NET39[27] NET39[28] NET39[29] NET39[30] 
+ NET39[31] NET39[32] NET39[33] NET39[34] NET39[35] NET39[36] NET39[37] 
+ NET39[38] NET39[39] NET39[40] NET39[41] NET39[42] NET39[43] NET39[44] 
+ NET39[45] NET39[46] NET39[47] NET39[48] NET39[49] NET39[50] NET39[51] 
+ NET39[52] NET39[53] NET39[54] NET39[55] NET39[56] NET39[57] NET39[58] 
+ NET39[59] NET39[60] NET39[61] NET39[62] NET39[63] WLPY_0UP[0] WLPYB_0UP[0] 
+ S1AHSF400W40_WLDV_64X1
XI3 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] PD_BUF PD_CVDDBUF VDDHD VDDI VSSI NET89[0] NET89[1] 
+ NET89[2] NET89[3] NET89[4] NET89[5] NET89[6] NET89[7] NET89[8] NET89[9] 
+ NET89[10] NET89[11] NET89[12] NET89[13] NET89[14] NET89[15] NET89[16] 
+ NET89[17] NET89[18] NET89[19] NET89[20] NET89[21] NET89[22] NET89[23] 
+ NET89[24] NET89[25] NET89[26] NET89[27] NET89[28] NET89[29] NET89[30] 
+ NET89[31] NET89[32] NET89[33] NET89[34] NET89[35] NET89[36] NET89[37] 
+ NET89[38] NET89[39] NET89[40] NET89[41] NET89[42] NET89[43] NET89[44] 
+ NET89[45] NET89[46] NET89[47] NET89[48] NET89[49] NET89[50] NET89[51] 
+ NET89[52] NET89[53] NET89[54] NET89[55] NET89[56] NET89[57] NET89[58] 
+ NET89[59] NET89[60] NET89[61] NET89[62] NET89[63] WLPY_3DN[0] WLPYB_3DN[0] 
+ S1AHSF400W40_WLDV_64X1
XI1 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] PD_BUF PD_CVDDBUF VDDHD VDDI VSSI NET49[0] NET49[1] 
+ NET49[2] NET49[3] NET49[4] NET49[5] NET49[6] NET49[7] NET49[8] NET49[9] 
+ NET49[10] NET49[11] NET49[12] NET49[13] NET49[14] NET49[15] NET49[16] 
+ NET49[17] NET49[18] NET49[19] NET49[20] NET49[21] NET49[22] NET49[23] 
+ NET49[24] NET49[25] NET49[26] NET49[27] NET49[28] NET49[29] NET49[30] 
+ NET49[31] NET49[32] NET49[33] NET49[34] NET49[35] NET49[36] NET49[37] 
+ NET49[38] NET49[39] NET49[40] NET49[41] NET49[42] NET49[43] NET49[44] 
+ NET49[45] NET49[46] NET49[47] NET49[48] NET49[49] NET49[50] NET49[51] 
+ NET49[52] NET49[53] NET49[54] NET49[55] NET49[56] NET49[57] NET49[58] 
+ NET49[59] NET49[60] NET49[61] NET49[62] NET49[63] WLPY_1DN[0] WLPYB_1DN[0] 
+ S1AHSF400W40_WLDV_64X1
XI0 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] PD_BUF PD_CVDDBUF VDDHD VDDI VSSI NET59[0] NET59[1] 
+ NET59[2] NET59[3] NET59[4] NET59[5] NET59[6] NET59[7] NET59[8] NET59[9] 
+ NET59[10] NET59[11] NET59[12] NET59[13] NET59[14] NET59[15] NET59[16] 
+ NET59[17] NET59[18] NET59[19] NET59[20] NET59[21] NET59[22] NET59[23] 
+ NET59[24] NET59[25] NET59[26] NET59[27] NET59[28] NET59[29] NET59[30] 
+ NET59[31] NET59[32] NET59[33] NET59[34] NET59[35] NET59[36] NET59[37] 
+ NET59[38] NET59[39] NET59[40] NET59[41] NET59[42] NET59[43] NET59[44] 
+ NET59[45] NET59[46] NET59[47] NET59[48] NET59[49] NET59[50] NET59[51] 
+ NET59[52] NET59[53] NET59[54] NET59[55] NET59[56] NET59[57] NET59[58] 
+ NET59[59] NET59[60] NET59[61] NET59[62] NET59[63] WLPY_1UP[0] WLPYB_1UP[0] 
+ S1AHSF400W40_WLDV_64X1
XWLDV_256X1_U DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] PD_BUF PD_CVDDBUF VDDHD VDDI VSSI NET79[0] 
+ NET79[1] NET79[2] NET79[3] NET79[4] NET79[5] NET79[6] NET79[7] NET79[8] 
+ NET79[9] NET79[10] NET79[11] NET79[12] NET79[13] NET79[14] NET79[15] 
+ NET79[16] NET79[17] NET79[18] NET79[19] NET79[20] NET79[21] NET79[22] 
+ NET79[23] NET79[24] NET79[25] NET79[26] NET79[27] NET79[28] NET79[29] 
+ NET79[30] NET79[31] NET79[32] NET79[33] NET79[34] NET79[35] NET79[36] 
+ NET79[37] NET79[38] NET79[39] NET79[40] NET79[41] NET79[42] NET79[43] 
+ NET79[44] NET79[45] NET79[46] NET79[47] NET79[48] NET79[49] NET79[50] 
+ NET79[51] NET79[52] NET79[53] NET79[54] NET79[55] NET79[56] NET79[57] 
+ NET79[58] NET79[59] NET79[60] NET79[61] NET79[62] NET79[63] WLPY_2UP[0] 
+ WLPYB_2UP[0] S1AHSF400W40_WLDV_64X1
XWLDV_256X1_D DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] PD_BUF PD_CVDDBUF VDDHD VDDI VSSI NET69[0] 
+ NET69[1] NET69[2] NET69[3] NET69[4] NET69[5] NET69[6] NET69[7] NET69[8] 
+ NET69[9] NET69[10] NET69[11] NET69[12] NET69[13] NET69[14] NET69[15] 
+ NET69[16] NET69[17] NET69[18] NET69[19] NET69[20] NET69[21] NET69[22] 
+ NET69[23] NET69[24] NET69[25] NET69[26] NET69[27] NET69[28] NET69[29] 
+ NET69[30] NET69[31] NET69[32] NET69[33] NET69[34] NET69[35] NET69[36] 
+ NET69[37] NET69[38] NET69[39] NET69[40] NET69[41] NET69[42] NET69[43] 
+ NET69[44] NET69[45] NET69[46] NET69[47] NET69[48] NET69[49] NET69[50] 
+ NET69[51] NET69[52] NET69[53] NET69[54] NET69[55] NET69[56] NET69[57] 
+ NET69[58] NET69[59] NET69[60] NET69[61] NET69[62] NET69[63] WLPY_2DN[0] 
+ WLPYB_2DN[0] S1AHSF400W40_WLDV_64X1
XI2 NET135 NET133 NET097[0] NET097[1] NET097[2] NET097[3] NET097[4] NET097[5] 
+ NET097[6] NET097[7] NET096[0] NET096[1] NET096[2] NET096[3] NET096[4] 
+ NET096[5] NET096[6] NET096[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] 
+ DEC_X3[2] DEC_X3[3] NET093[0] NET093[1] NET093[2] NET093[3] NET093[4] 
+ NET093[5] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] 
+ DEC_Y[7] NET131[0] NET131[1] NET131[2] NET131[3] NET131[4] NET131[5] 
+ NET131[6] NET131[7] NET136[0] NET136[1] NET136[2] NET136[3] NET136[4] 
+ NET136[5] NET136[6] NET136[7] PD_BUF PD_CVDDBUF NET137 RW_RE NET132 VDDHD 
+ VDDI VSSI NET134 WLPY_1DN[0] WLPY_1DN[1] WLPY_1DN[2] WLPY_1DN[3] WLPY_1UP[0] 
+ WLPY_1UP[1] WLPY_1UP[2] WLPY_1UP[3] WLP_SAE NET010 YL[0] NET122[0] NET122[1] 
+ S1AHSF400W40_LCTRL_F_M4
XLCTRL_S_M4 NET31 NET29 NET0122[0] NET0122[1] NET0122[2] NET0122[3] NET0122[4] 
+ NET0122[5] NET0122[6] NET0122[7] NET0121[0] NET0121[1] NET0121[2] NET0121[3] 
+ NET0121[4] NET0121[5] NET0121[6] NET0121[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[4] DEC_X3[5] NET0118[0] NET0118[1] NET0118[2] NET0118[3] 
+ NET0118[4] NET0118[5] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] NET27[0] NET27[1] NET27[2] NET27[3] NET27[4] NET27[5] 
+ NET27[6] NET27[7] NET32[0] NET32[1] NET32[2] NET32[3] NET32[4] NET32[5] 
+ NET32[6] NET32[7] PD_BUF PD_CVDDBUF NET33 RW_RE NET28 VDDHD VDDI VSSI NET30 
+ WLPY_2DN[0] WLPY_2DN[1] WLPY_2DN[2] WLPY_2DN[3] WLPY_2UP[0] WLPY_2UP[1] 
+ WLPY_2UP[2] WLPY_2UP[3] WLP_SAE NET0119 YL[0] NET18[0] NET18[1] S1AHSF400W40_LCTRL_F_M4
XXDRV_STRP_1D VDDHD VDDI VSSI WLPY_1DN[0] WLPYB_1DN[0] S1AHSF400W40_XDRV_STRAP
XI7 VDDHD VDDI VSSI WLPY_2UP[0] WLPYB_2UP[0] S1AHSF400W40_XDRV_STRAP
XI6 VDDHD VDDI VSSI WLPY_2DN[0] WLPYB_2DN[0] S1AHSF400W40_XDRV_STRAP
XXDRV_STRAP_1U<0> VDDHD VDDI VSSI WLPY_1UP[0] WLPYB_1UP[0] S1AHSF400W40_XDRV_STRAP
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    WLDV_256X1
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_WLDV_256X1 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] PD_BUF PD_CVDDBUF VDDHD VDDI VSSI WL[0] WL[1] 
+ WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] 
+ WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] 
+ WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] 
+ WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] 
+ WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] 
+ WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] 
+ WL[69] WL[70] WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] 
+ WL[80] WL[81] WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] 
+ WL[91] WL[92] WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] 
+ WL[101] WL[102] WL[103] WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] 
+ WL[110] WL[111] WL[112] WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] 
+ WL[119] WL[120] WL[121] WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] 
+ WL[128] WL[129] WL[130] WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] 
+ WL[137] WL[138] WL[139] WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] 
+ WL[146] WL[147] WL[148] WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] 
+ WL[155] WL[156] WL[157] WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] 
+ WL[164] WL[165] WL[166] WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] 
+ WL[173] WL[174] WL[175] WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] 
+ WL[182] WL[183] WL[184] WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] 
+ WL[191] WL[192] WL[193] WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] 
+ WL[200] WL[201] WL[202] WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] 
+ WL[209] WL[210] WL[211] WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] 
+ WL[218] WL[219] WL[220] WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] 
+ WL[227] WL[228] WL[229] WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] 
+ WL[236] WL[237] WL[238] WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] 
+ WL[245] WL[246] WL[247] WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] 
+ WL[254] WL[255] WLPY[0] WLPY[1] WLPY[2] WLPY[3] WLPYB[0] WLPYB[1] WLPYB[2] 
+ WLPYB[3]
*.PININFO DEC_X0[0]:I DEC_X0[1]:I DEC_X0[2]:I DEC_X0[3]:I DEC_X0[4]:I 
*.PININFO DEC_X0[5]:I DEC_X0[6]:I DEC_X0[7]:I DEC_X1[0]:I DEC_X1[1]:I 
*.PININFO DEC_X1[2]:I DEC_X1[3]:I DEC_X1[4]:I DEC_X1[5]:I DEC_X1[6]:I 
*.PININFO DEC_X1[7]:I PD_BUF:I PD_CVDDBUF:I WLPY[0]:I WLPY[1]:I WLPY[2]:I 
*.PININFO WLPY[3]:I WLPYB[0]:I WLPYB[1]:I WLPYB[2]:I WLPYB[3]:I WL[0]:O 
*.PININFO WL[1]:O WL[2]:O WL[3]:O WL[4]:O WL[5]:O WL[6]:O WL[7]:O WL[8]:O 
*.PININFO WL[9]:O WL[10]:O WL[11]:O WL[12]:O WL[13]:O WL[14]:O WL[15]:O 
*.PININFO WL[16]:O WL[17]:O WL[18]:O WL[19]:O WL[20]:O WL[21]:O WL[22]:O 
*.PININFO WL[23]:O WL[24]:O WL[25]:O WL[26]:O WL[27]:O WL[28]:O WL[29]:O 
*.PININFO WL[30]:O WL[31]:O WL[32]:O WL[33]:O WL[34]:O WL[35]:O WL[36]:O 
*.PININFO WL[37]:O WL[38]:O WL[39]:O WL[40]:O WL[41]:O WL[42]:O WL[43]:O 
*.PININFO WL[44]:O WL[45]:O WL[46]:O WL[47]:O WL[48]:O WL[49]:O WL[50]:O 
*.PININFO WL[51]:O WL[52]:O WL[53]:O WL[54]:O WL[55]:O WL[56]:O WL[57]:O 
*.PININFO WL[58]:O WL[59]:O WL[60]:O WL[61]:O WL[62]:O WL[63]:O WL[64]:O 
*.PININFO WL[65]:O WL[66]:O WL[67]:O WL[68]:O WL[69]:O WL[70]:O WL[71]:O 
*.PININFO WL[72]:O WL[73]:O WL[74]:O WL[75]:O WL[76]:O WL[77]:O WL[78]:O 
*.PININFO WL[79]:O WL[80]:O WL[81]:O WL[82]:O WL[83]:O WL[84]:O WL[85]:O 
*.PININFO WL[86]:O WL[87]:O WL[88]:O WL[89]:O WL[90]:O WL[91]:O WL[92]:O 
*.PININFO WL[93]:O WL[94]:O WL[95]:O WL[96]:O WL[97]:O WL[98]:O WL[99]:O 
*.PININFO WL[100]:O WL[101]:O WL[102]:O WL[103]:O WL[104]:O WL[105]:O 
*.PININFO WL[106]:O WL[107]:O WL[108]:O WL[109]:O WL[110]:O WL[111]:O 
*.PININFO WL[112]:O WL[113]:O WL[114]:O WL[115]:O WL[116]:O WL[117]:O 
*.PININFO WL[118]:O WL[119]:O WL[120]:O WL[121]:O WL[122]:O WL[123]:O 
*.PININFO WL[124]:O WL[125]:O WL[126]:O WL[127]:O WL[128]:O WL[129]:O 
*.PININFO WL[130]:O WL[131]:O WL[132]:O WL[133]:O WL[134]:O WL[135]:O 
*.PININFO WL[136]:O WL[137]:O WL[138]:O WL[139]:O WL[140]:O WL[141]:O 
*.PININFO WL[142]:O WL[143]:O WL[144]:O WL[145]:O WL[146]:O WL[147]:O 
*.PININFO WL[148]:O WL[149]:O WL[150]:O WL[151]:O WL[152]:O WL[153]:O 
*.PININFO WL[154]:O WL[155]:O WL[156]:O WL[157]:O WL[158]:O WL[159]:O 
*.PININFO WL[160]:O WL[161]:O WL[162]:O WL[163]:O WL[164]:O WL[165]:O 
*.PININFO WL[166]:O WL[167]:O WL[168]:O WL[169]:O WL[170]:O WL[171]:O 
*.PININFO WL[172]:O WL[173]:O WL[174]:O WL[175]:O WL[176]:O WL[177]:O 
*.PININFO WL[178]:O WL[179]:O WL[180]:O WL[181]:O WL[182]:O WL[183]:O 
*.PININFO WL[184]:O WL[185]:O WL[186]:O WL[187]:O WL[188]:O WL[189]:O 
*.PININFO WL[190]:O WL[191]:O WL[192]:O WL[193]:O WL[194]:O WL[195]:O 
*.PININFO WL[196]:O WL[197]:O WL[198]:O WL[199]:O WL[200]:O WL[201]:O 
*.PININFO WL[202]:O WL[203]:O WL[204]:O WL[205]:O WL[206]:O WL[207]:O 
*.PININFO WL[208]:O WL[209]:O WL[210]:O WL[211]:O WL[212]:O WL[213]:O 
*.PININFO WL[214]:O WL[215]:O WL[216]:O WL[217]:O WL[218]:O WL[219]:O 
*.PININFO WL[220]:O WL[221]:O WL[222]:O WL[223]:O WL[224]:O WL[225]:O 
*.PININFO WL[226]:O WL[227]:O WL[228]:O WL[229]:O WL[230]:O WL[231]:O 
*.PININFO WL[232]:O WL[233]:O WL[234]:O WL[235]:O WL[236]:O WL[237]:O 
*.PININFO WL[238]:O WL[239]:O WL[240]:O WL[241]:O WL[242]:O WL[243]:O 
*.PININFO WL[244]:O WL[245]:O WL[246]:O WL[247]:O WL[248]:O WL[249]:O 
*.PININFO WL[250]:O WL[251]:O WL[252]:O WL[253]:O WL[254]:O WL[255]:O VDDHD:B 
*.PININFO VDDI:B VSSI:B
XWLDV_2X1<16> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[0] NET17[0] 
+ NET17[1] NET17[2] NET17[3] NET16[0] NET16[1] NET16[2] NET16[3] NET16[4] 
+ NET16[5] NET16[6] NET16[7] NET15[0] NET15[1] NET15[2] NET15[3] NET15[4] 
+ NET15[5] NET15[6] NET15[7] PD_BUF PD_CVDDBUF NET14[0] VDDHD VDDI VSSI WL[64] 
+ WL[65] WL[66] WL[67] WLPY[1] WLPYB[1] NET13[0] NET12[0] NET11[0] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<17> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] NET17[4] 
+ NET17[5] NET17[6] NET17[7] NET16[8] NET16[9] NET16[10] NET16[11] NET16[12] 
+ NET16[13] NET16[14] NET16[15] NET15[8] NET15[9] NET15[10] NET15[11] 
+ NET15[12] NET15[13] NET15[14] NET15[15] PD_BUF PD_CVDDBUF NET14[1] VDDHD 
+ VDDI VSSI WL[68] WL[69] WL[70] WL[71] WLPY[1] WLPYB[1] NET13[1] NET12[1] 
+ NET11[1] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<18> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[1] NET17[8] 
+ NET17[9] NET17[10] NET17[11] NET16[16] NET16[17] NET16[18] NET16[19] 
+ NET16[20] NET16[21] NET16[22] NET16[23] NET15[16] NET15[17] NET15[18] 
+ NET15[19] NET15[20] NET15[21] NET15[22] NET15[23] PD_BUF PD_CVDDBUF NET14[2] 
+ VDDHD VDDI VSSI WL[72] WL[73] WL[74] WL[75] WLPY[1] WLPYB[1] NET13[2] 
+ NET12[2] NET11[2] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<19> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] NET17[12] 
+ NET17[13] NET17[14] NET17[15] NET16[24] NET16[25] NET16[26] NET16[27] 
+ NET16[28] NET16[29] NET16[30] NET16[31] NET15[24] NET15[25] NET15[26] 
+ NET15[27] NET15[28] NET15[29] NET15[30] NET15[31] PD_BUF PD_CVDDBUF NET14[3] 
+ VDDHD VDDI VSSI WL[76] WL[77] WL[78] WL[79] WLPY[1] WLPYB[1] NET13[3] 
+ NET12[3] NET11[3] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<20> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[2] NET17[16] 
+ NET17[17] NET17[18] NET17[19] NET16[32] NET16[33] NET16[34] NET16[35] 
+ NET16[36] NET16[37] NET16[38] NET16[39] NET15[32] NET15[33] NET15[34] 
+ NET15[35] NET15[36] NET15[37] NET15[38] NET15[39] PD_BUF PD_CVDDBUF NET14[4] 
+ VDDHD VDDI VSSI WL[80] WL[81] WL[82] WL[83] WLPY[1] WLPYB[1] NET13[4] 
+ NET12[4] NET11[4] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<21> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] NET17[20] 
+ NET17[21] NET17[22] NET17[23] NET16[40] NET16[41] NET16[42] NET16[43] 
+ NET16[44] NET16[45] NET16[46] NET16[47] NET15[40] NET15[41] NET15[42] 
+ NET15[43] NET15[44] NET15[45] NET15[46] NET15[47] PD_BUF PD_CVDDBUF NET14[5] 
+ VDDHD VDDI VSSI WL[84] WL[85] WL[86] WL[87] WLPY[1] WLPYB[1] NET13[5] 
+ NET12[5] NET11[5] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<22> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[3] NET17[24] 
+ NET17[25] NET17[26] NET17[27] NET16[48] NET16[49] NET16[50] NET16[51] 
+ NET16[52] NET16[53] NET16[54] NET16[55] NET15[48] NET15[49] NET15[50] 
+ NET15[51] NET15[52] NET15[53] NET15[54] NET15[55] PD_BUF PD_CVDDBUF NET14[6] 
+ VDDHD VDDI VSSI WL[88] WL[89] WL[90] WL[91] WLPY[1] WLPYB[1] NET13[6] 
+ NET12[6] NET11[6] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<23> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] NET17[28] 
+ NET17[29] NET17[30] NET17[31] NET16[56] NET16[57] NET16[58] NET16[59] 
+ NET16[60] NET16[61] NET16[62] NET16[63] NET15[56] NET15[57] NET15[58] 
+ NET15[59] NET15[60] NET15[61] NET15[62] NET15[63] PD_BUF PD_CVDDBUF NET14[7] 
+ VDDHD VDDI VSSI WL[92] WL[93] WL[94] WL[95] WLPY[1] WLPYB[1] NET13[7] 
+ NET12[7] NET11[7] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<24> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[4] NET17[32] 
+ NET17[33] NET17[34] NET17[35] NET16[64] NET16[65] NET16[66] NET16[67] 
+ NET16[68] NET16[69] NET16[70] NET16[71] NET15[64] NET15[65] NET15[66] 
+ NET15[67] NET15[68] NET15[69] NET15[70] NET15[71] PD_BUF PD_CVDDBUF NET14[8] 
+ VDDHD VDDI VSSI WL[96] WL[97] WL[98] WL[99] WLPY[1] WLPYB[1] NET13[8] 
+ NET12[8] NET11[8] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<25> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] NET17[36] 
+ NET17[37] NET17[38] NET17[39] NET16[72] NET16[73] NET16[74] NET16[75] 
+ NET16[76] NET16[77] NET16[78] NET16[79] NET15[72] NET15[73] NET15[74] 
+ NET15[75] NET15[76] NET15[77] NET15[78] NET15[79] PD_BUF PD_CVDDBUF NET14[9] 
+ VDDHD VDDI VSSI WL[100] WL[101] WL[102] WL[103] WLPY[1] WLPYB[1] NET13[9] 
+ NET12[9] NET11[9] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<26> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[5] NET17[40] 
+ NET17[41] NET17[42] NET17[43] NET16[80] NET16[81] NET16[82] NET16[83] 
+ NET16[84] NET16[85] NET16[86] NET16[87] NET15[80] NET15[81] NET15[82] 
+ NET15[83] NET15[84] NET15[85] NET15[86] NET15[87] PD_BUF PD_CVDDBUF 
+ NET14[10] VDDHD VDDI VSSI WL[104] WL[105] WL[106] WL[107] WLPY[1] WLPYB[1] 
+ NET13[10] NET12[10] NET11[10] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<27> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] NET17[44] 
+ NET17[45] NET17[46] NET17[47] NET16[88] NET16[89] NET16[90] NET16[91] 
+ NET16[92] NET16[93] NET16[94] NET16[95] NET15[88] NET15[89] NET15[90] 
+ NET15[91] NET15[92] NET15[93] NET15[94] NET15[95] PD_BUF PD_CVDDBUF 
+ NET14[11] VDDHD VDDI VSSI WL[108] WL[109] WL[110] WL[111] WLPY[1] WLPYB[1] 
+ NET13[11] NET12[11] NET11[11] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<28> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[6] NET17[48] 
+ NET17[49] NET17[50] NET17[51] NET16[96] NET16[97] NET16[98] NET16[99] 
+ NET16[100] NET16[101] NET16[102] NET16[103] NET15[96] NET15[97] NET15[98] 
+ NET15[99] NET15[100] NET15[101] NET15[102] NET15[103] PD_BUF PD_CVDDBUF 
+ NET14[12] VDDHD VDDI VSSI WL[112] WL[113] WL[114] WL[115] WLPY[1] WLPYB[1] 
+ NET13[12] NET12[12] NET11[12] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<29> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] NET17[52] 
+ NET17[53] NET17[54] NET17[55] NET16[104] NET16[105] NET16[106] NET16[107] 
+ NET16[108] NET16[109] NET16[110] NET16[111] NET15[104] NET15[105] NET15[106] 
+ NET15[107] NET15[108] NET15[109] NET15[110] NET15[111] PD_BUF PD_CVDDBUF 
+ NET14[13] VDDHD VDDI VSSI WL[116] WL[117] WL[118] WL[119] WLPY[1] WLPYB[1] 
+ NET13[13] NET12[13] NET11[13] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<30> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[7] NET17[56] 
+ NET17[57] NET17[58] NET17[59] NET16[112] NET16[113] NET16[114] NET16[115] 
+ NET16[116] NET16[117] NET16[118] NET16[119] NET15[112] NET15[113] NET15[114] 
+ NET15[115] NET15[116] NET15[117] NET15[118] NET15[119] PD_BUF PD_CVDDBUF 
+ NET14[14] VDDHD VDDI VSSI WL[120] WL[121] WL[122] WL[123] WLPY[1] WLPYB[1] 
+ NET13[14] NET12[14] NET11[14] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<31> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] NET17[60] 
+ NET17[61] NET17[62] NET17[63] NET16[120] NET16[121] NET16[122] NET16[123] 
+ NET16[124] NET16[125] NET16[126] NET16[127] NET15[120] NET15[121] NET15[122] 
+ NET15[123] NET15[124] NET15[125] NET15[126] NET15[127] PD_BUF PD_CVDDBUF 
+ NET14[15] VDDHD VDDI VSSI WL[124] WL[125] WL[126] WL[127] WLPY[1] WLPYB[1] 
+ NET13[15] NET12[15] NET11[15] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<32> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[0] NET34[0] 
+ NET34[1] NET34[2] NET34[3] NET33[0] NET33[1] NET33[2] NET33[3] NET33[4] 
+ NET33[5] NET33[6] NET33[7] NET32[0] NET32[1] NET32[2] NET32[3] NET32[4] 
+ NET32[5] NET32[6] NET32[7] PD_BUF PD_CVDDBUF NET31[0] VDDHD VDDI VSSI 
+ WL[128] WL[129] WL[130] WL[131] WLPY[2] WLPYB[2] NET30[0] NET29[0] NET28[0] 
+ S1AHSF400W40_WLDV_2X1
XWLDV_2X1<33> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] NET34[4] 
+ NET34[5] NET34[6] NET34[7] NET33[8] NET33[9] NET33[10] NET33[11] NET33[12] 
+ NET33[13] NET33[14] NET33[15] NET32[8] NET32[9] NET32[10] NET32[11] 
+ NET32[12] NET32[13] NET32[14] NET32[15] PD_BUF PD_CVDDBUF NET31[1] VDDHD 
+ VDDI VSSI WL[132] WL[133] WL[134] WL[135] WLPY[2] WLPYB[2] NET30[1] NET29[1] 
+ NET28[1] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<34> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[1] NET34[8] 
+ NET34[9] NET34[10] NET34[11] NET33[16] NET33[17] NET33[18] NET33[19] 
+ NET33[20] NET33[21] NET33[22] NET33[23] NET32[16] NET32[17] NET32[18] 
+ NET32[19] NET32[20] NET32[21] NET32[22] NET32[23] PD_BUF PD_CVDDBUF NET31[2] 
+ VDDHD VDDI VSSI WL[136] WL[137] WL[138] WL[139] WLPY[2] WLPYB[2] NET30[2] 
+ NET29[2] NET28[2] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<35> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] NET34[12] 
+ NET34[13] NET34[14] NET34[15] NET33[24] NET33[25] NET33[26] NET33[27] 
+ NET33[28] NET33[29] NET33[30] NET33[31] NET32[24] NET32[25] NET32[26] 
+ NET32[27] NET32[28] NET32[29] NET32[30] NET32[31] PD_BUF PD_CVDDBUF NET31[3] 
+ VDDHD VDDI VSSI WL[140] WL[141] WL[142] WL[143] WLPY[2] WLPYB[2] NET30[3] 
+ NET29[3] NET28[3] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<36> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[2] NET34[16] 
+ NET34[17] NET34[18] NET34[19] NET33[32] NET33[33] NET33[34] NET33[35] 
+ NET33[36] NET33[37] NET33[38] NET33[39] NET32[32] NET32[33] NET32[34] 
+ NET32[35] NET32[36] NET32[37] NET32[38] NET32[39] PD_BUF PD_CVDDBUF NET31[4] 
+ VDDHD VDDI VSSI WL[144] WL[145] WL[146] WL[147] WLPY[2] WLPYB[2] NET30[4] 
+ NET29[4] NET28[4] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<37> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] NET34[20] 
+ NET34[21] NET34[22] NET34[23] NET33[40] NET33[41] NET33[42] NET33[43] 
+ NET33[44] NET33[45] NET33[46] NET33[47] NET32[40] NET32[41] NET32[42] 
+ NET32[43] NET32[44] NET32[45] NET32[46] NET32[47] PD_BUF PD_CVDDBUF NET31[5] 
+ VDDHD VDDI VSSI WL[148] WL[149] WL[150] WL[151] WLPY[2] WLPYB[2] NET30[5] 
+ NET29[5] NET28[5] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<38> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[3] NET34[24] 
+ NET34[25] NET34[26] NET34[27] NET33[48] NET33[49] NET33[50] NET33[51] 
+ NET33[52] NET33[53] NET33[54] NET33[55] NET32[48] NET32[49] NET32[50] 
+ NET32[51] NET32[52] NET32[53] NET32[54] NET32[55] PD_BUF PD_CVDDBUF NET31[6] 
+ VDDHD VDDI VSSI WL[152] WL[153] WL[154] WL[155] WLPY[2] WLPYB[2] NET30[6] 
+ NET29[6] NET28[6] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<39> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] NET34[28] 
+ NET34[29] NET34[30] NET34[31] NET33[56] NET33[57] NET33[58] NET33[59] 
+ NET33[60] NET33[61] NET33[62] NET33[63] NET32[56] NET32[57] NET32[58] 
+ NET32[59] NET32[60] NET32[61] NET32[62] NET32[63] PD_BUF PD_CVDDBUF NET31[7] 
+ VDDHD VDDI VSSI WL[156] WL[157] WL[158] WL[159] WLPY[2] WLPYB[2] NET30[7] 
+ NET29[7] NET28[7] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<40> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[4] NET34[32] 
+ NET34[33] NET34[34] NET34[35] NET33[64] NET33[65] NET33[66] NET33[67] 
+ NET33[68] NET33[69] NET33[70] NET33[71] NET32[64] NET32[65] NET32[66] 
+ NET32[67] NET32[68] NET32[69] NET32[70] NET32[71] PD_BUF PD_CVDDBUF NET31[8] 
+ VDDHD VDDI VSSI WL[160] WL[161] WL[162] WL[163] WLPY[2] WLPYB[2] NET30[8] 
+ NET29[8] NET28[8] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<41> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] NET34[36] 
+ NET34[37] NET34[38] NET34[39] NET33[72] NET33[73] NET33[74] NET33[75] 
+ NET33[76] NET33[77] NET33[78] NET33[79] NET32[72] NET32[73] NET32[74] 
+ NET32[75] NET32[76] NET32[77] NET32[78] NET32[79] PD_BUF PD_CVDDBUF NET31[9] 
+ VDDHD VDDI VSSI WL[164] WL[165] WL[166] WL[167] WLPY[2] WLPYB[2] NET30[9] 
+ NET29[9] NET28[9] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<42> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[5] NET34[40] 
+ NET34[41] NET34[42] NET34[43] NET33[80] NET33[81] NET33[82] NET33[83] 
+ NET33[84] NET33[85] NET33[86] NET33[87] NET32[80] NET32[81] NET32[82] 
+ NET32[83] NET32[84] NET32[85] NET32[86] NET32[87] PD_BUF PD_CVDDBUF 
+ NET31[10] VDDHD VDDI VSSI WL[168] WL[169] WL[170] WL[171] WLPY[2] WLPYB[2] 
+ NET30[10] NET29[10] NET28[10] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<43> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] NET34[44] 
+ NET34[45] NET34[46] NET34[47] NET33[88] NET33[89] NET33[90] NET33[91] 
+ NET33[92] NET33[93] NET33[94] NET33[95] NET32[88] NET32[89] NET32[90] 
+ NET32[91] NET32[92] NET32[93] NET32[94] NET32[95] PD_BUF PD_CVDDBUF 
+ NET31[11] VDDHD VDDI VSSI WL[172] WL[173] WL[174] WL[175] WLPY[2] WLPYB[2] 
+ NET30[11] NET29[11] NET28[11] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<44> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[6] NET34[48] 
+ NET34[49] NET34[50] NET34[51] NET33[96] NET33[97] NET33[98] NET33[99] 
+ NET33[100] NET33[101] NET33[102] NET33[103] NET32[96] NET32[97] NET32[98] 
+ NET32[99] NET32[100] NET32[101] NET32[102] NET32[103] PD_BUF PD_CVDDBUF 
+ NET31[12] VDDHD VDDI VSSI WL[176] WL[177] WL[178] WL[179] WLPY[2] WLPYB[2] 
+ NET30[12] NET29[12] NET28[12] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<45> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] NET34[52] 
+ NET34[53] NET34[54] NET34[55] NET33[104] NET33[105] NET33[106] NET33[107] 
+ NET33[108] NET33[109] NET33[110] NET33[111] NET32[104] NET32[105] NET32[106] 
+ NET32[107] NET32[108] NET32[109] NET32[110] NET32[111] PD_BUF PD_CVDDBUF 
+ NET31[13] VDDHD VDDI VSSI WL[180] WL[181] WL[182] WL[183] WLPY[2] WLPYB[2] 
+ NET30[13] NET29[13] NET28[13] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<46> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[7] NET34[56] 
+ NET34[57] NET34[58] NET34[59] NET33[112] NET33[113] NET33[114] NET33[115] 
+ NET33[116] NET33[117] NET33[118] NET33[119] NET32[112] NET32[113] NET32[114] 
+ NET32[115] NET32[116] NET32[117] NET32[118] NET32[119] PD_BUF PD_CVDDBUF 
+ NET31[14] VDDHD VDDI VSSI WL[184] WL[185] WL[186] WL[187] WLPY[2] WLPYB[2] 
+ NET30[14] NET29[14] NET28[14] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<47> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] NET34[60] 
+ NET34[61] NET34[62] NET34[63] NET33[120] NET33[121] NET33[122] NET33[123] 
+ NET33[124] NET33[125] NET33[126] NET33[127] NET32[120] NET32[121] NET32[122] 
+ NET32[123] NET32[124] NET32[125] NET32[126] NET32[127] PD_BUF PD_CVDDBUF 
+ NET31[15] VDDHD VDDI VSSI WL[188] WL[189] WL[190] WL[191] WLPY[2] WLPYB[2] 
+ NET30[15] NET29[15] NET28[15] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<0> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[0] NET51[0] 
+ NET51[1] NET51[2] NET51[3] NET50[0] NET50[1] NET50[2] NET50[3] NET50[4] 
+ NET50[5] NET50[6] NET50[7] NET49[0] NET49[1] NET49[2] NET49[3] NET49[4] 
+ NET49[5] NET49[6] NET49[7] PD_BUF PD_CVDDBUF NET48[0] VDDHD VDDI VSSI WL[0] 
+ WL[1] WL[2] WL[3] WLPY[0] WLPYB[0] NET47[0] NET46[0] NET45[0] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<1> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] NET51[4] 
+ NET51[5] NET51[6] NET51[7] NET50[8] NET50[9] NET50[10] NET50[11] NET50[12] 
+ NET50[13] NET50[14] NET50[15] NET49[8] NET49[9] NET49[10] NET49[11] 
+ NET49[12] NET49[13] NET49[14] NET49[15] PD_BUF PD_CVDDBUF NET48[1] VDDHD 
+ VDDI VSSI WL[4] WL[5] WL[6] WL[7] WLPY[0] WLPYB[0] NET47[1] NET46[1] 
+ NET45[1] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<2> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[1] NET51[8] 
+ NET51[9] NET51[10] NET51[11] NET50[16] NET50[17] NET50[18] NET50[19] 
+ NET50[20] NET50[21] NET50[22] NET50[23] NET49[16] NET49[17] NET49[18] 
+ NET49[19] NET49[20] NET49[21] NET49[22] NET49[23] PD_BUF PD_CVDDBUF NET48[2] 
+ VDDHD VDDI VSSI WL[8] WL[9] WL[10] WL[11] WLPY[0] WLPYB[0] NET47[2] NET46[2] 
+ NET45[2] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<3> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] NET51[12] 
+ NET51[13] NET51[14] NET51[15] NET50[24] NET50[25] NET50[26] NET50[27] 
+ NET50[28] NET50[29] NET50[30] NET50[31] NET49[24] NET49[25] NET49[26] 
+ NET49[27] NET49[28] NET49[29] NET49[30] NET49[31] PD_BUF PD_CVDDBUF NET48[3] 
+ VDDHD VDDI VSSI WL[12] WL[13] WL[14] WL[15] WLPY[0] WLPYB[0] NET47[3] 
+ NET46[3] NET45[3] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<4> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[2] NET51[16] 
+ NET51[17] NET51[18] NET51[19] NET50[32] NET50[33] NET50[34] NET50[35] 
+ NET50[36] NET50[37] NET50[38] NET50[39] NET49[32] NET49[33] NET49[34] 
+ NET49[35] NET49[36] NET49[37] NET49[38] NET49[39] PD_BUF PD_CVDDBUF NET48[4] 
+ VDDHD VDDI VSSI WL[16] WL[17] WL[18] WL[19] WLPY[0] WLPYB[0] NET47[4] 
+ NET46[4] NET45[4] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<5> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] NET51[20] 
+ NET51[21] NET51[22] NET51[23] NET50[40] NET50[41] NET50[42] NET50[43] 
+ NET50[44] NET50[45] NET50[46] NET50[47] NET49[40] NET49[41] NET49[42] 
+ NET49[43] NET49[44] NET49[45] NET49[46] NET49[47] PD_BUF PD_CVDDBUF NET48[5] 
+ VDDHD VDDI VSSI WL[20] WL[21] WL[22] WL[23] WLPY[0] WLPYB[0] NET47[5] 
+ NET46[5] NET45[5] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<6> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[3] NET51[24] 
+ NET51[25] NET51[26] NET51[27] NET50[48] NET50[49] NET50[50] NET50[51] 
+ NET50[52] NET50[53] NET50[54] NET50[55] NET49[48] NET49[49] NET49[50] 
+ NET49[51] NET49[52] NET49[53] NET49[54] NET49[55] PD_BUF PD_CVDDBUF NET48[6] 
+ VDDHD VDDI VSSI WL[24] WL[25] WL[26] WL[27] WLPY[0] WLPYB[0] NET47[6] 
+ NET46[6] NET45[6] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<7> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] NET51[28] 
+ NET51[29] NET51[30] NET51[31] NET50[56] NET50[57] NET50[58] NET50[59] 
+ NET50[60] NET50[61] NET50[62] NET50[63] NET49[56] NET49[57] NET49[58] 
+ NET49[59] NET49[60] NET49[61] NET49[62] NET49[63] PD_BUF PD_CVDDBUF NET48[7] 
+ VDDHD VDDI VSSI WL[28] WL[29] WL[30] WL[31] WLPY[0] WLPYB[0] NET47[7] 
+ NET46[7] NET45[7] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<8> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[4] NET51[32] 
+ NET51[33] NET51[34] NET51[35] NET50[64] NET50[65] NET50[66] NET50[67] 
+ NET50[68] NET50[69] NET50[70] NET50[71] NET49[64] NET49[65] NET49[66] 
+ NET49[67] NET49[68] NET49[69] NET49[70] NET49[71] PD_BUF PD_CVDDBUF NET48[8] 
+ VDDHD VDDI VSSI WL[32] WL[33] WL[34] WL[35] WLPY[0] WLPYB[0] NET47[8] 
+ NET46[8] NET45[8] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<9> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] NET51[36] 
+ NET51[37] NET51[38] NET51[39] NET50[72] NET50[73] NET50[74] NET50[75] 
+ NET50[76] NET50[77] NET50[78] NET50[79] NET49[72] NET49[73] NET49[74] 
+ NET49[75] NET49[76] NET49[77] NET49[78] NET49[79] PD_BUF PD_CVDDBUF NET48[9] 
+ VDDHD VDDI VSSI WL[36] WL[37] WL[38] WL[39] WLPY[0] WLPYB[0] NET47[9] 
+ NET46[9] NET45[9] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<10> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[5] NET51[40] 
+ NET51[41] NET51[42] NET51[43] NET50[80] NET50[81] NET50[82] NET50[83] 
+ NET50[84] NET50[85] NET50[86] NET50[87] NET49[80] NET49[81] NET49[82] 
+ NET49[83] NET49[84] NET49[85] NET49[86] NET49[87] PD_BUF PD_CVDDBUF 
+ NET48[10] VDDHD VDDI VSSI WL[40] WL[41] WL[42] WL[43] WLPY[0] WLPYB[0] 
+ NET47[10] NET46[10] NET45[10] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<11> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] NET51[44] 
+ NET51[45] NET51[46] NET51[47] NET50[88] NET50[89] NET50[90] NET50[91] 
+ NET50[92] NET50[93] NET50[94] NET50[95] NET49[88] NET49[89] NET49[90] 
+ NET49[91] NET49[92] NET49[93] NET49[94] NET49[95] PD_BUF PD_CVDDBUF 
+ NET48[11] VDDHD VDDI VSSI WL[44] WL[45] WL[46] WL[47] WLPY[0] WLPYB[0] 
+ NET47[11] NET46[11] NET45[11] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<12> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[6] NET51[48] 
+ NET51[49] NET51[50] NET51[51] NET50[96] NET50[97] NET50[98] NET50[99] 
+ NET50[100] NET50[101] NET50[102] NET50[103] NET49[96] NET49[97] NET49[98] 
+ NET49[99] NET49[100] NET49[101] NET49[102] NET49[103] PD_BUF PD_CVDDBUF 
+ NET48[12] VDDHD VDDI VSSI WL[48] WL[49] WL[50] WL[51] WLPY[0] WLPYB[0] 
+ NET47[12] NET46[12] NET45[12] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<13> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] NET51[52] 
+ NET51[53] NET51[54] NET51[55] NET50[104] NET50[105] NET50[106] NET50[107] 
+ NET50[108] NET50[109] NET50[110] NET50[111] NET49[104] NET49[105] NET49[106] 
+ NET49[107] NET49[108] NET49[109] NET49[110] NET49[111] PD_BUF PD_CVDDBUF 
+ NET48[13] VDDHD VDDI VSSI WL[52] WL[53] WL[54] WL[55] WLPY[0] WLPYB[0] 
+ NET47[13] NET46[13] NET45[13] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<14> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[7] NET51[56] 
+ NET51[57] NET51[58] NET51[59] NET50[112] NET50[113] NET50[114] NET50[115] 
+ NET50[116] NET50[117] NET50[118] NET50[119] NET49[112] NET49[113] NET49[114] 
+ NET49[115] NET49[116] NET49[117] NET49[118] NET49[119] PD_BUF PD_CVDDBUF 
+ NET48[14] VDDHD VDDI VSSI WL[56] WL[57] WL[58] WL[59] WLPY[0] WLPYB[0] 
+ NET47[14] NET46[14] NET45[14] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<15> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] NET51[60] 
+ NET51[61] NET51[62] NET51[63] NET50[120] NET50[121] NET50[122] NET50[123] 
+ NET50[124] NET50[125] NET50[126] NET50[127] NET49[120] NET49[121] NET49[122] 
+ NET49[123] NET49[124] NET49[125] NET49[126] NET49[127] PD_BUF PD_CVDDBUF 
+ NET48[15] VDDHD VDDI VSSI WL[60] WL[61] WL[62] WL[63] WLPY[0] WLPYB[0] 
+ NET47[15] NET46[15] NET45[15] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<48> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[0] NET68[0] 
+ NET68[1] NET68[2] NET68[3] NET67[0] NET67[1] NET67[2] NET67[3] NET67[4] 
+ NET67[5] NET67[6] NET67[7] NET66[0] NET66[1] NET66[2] NET66[3] NET66[4] 
+ NET66[5] NET66[6] NET66[7] PD_BUF PD_CVDDBUF NET65[0] VDDHD VDDI VSSI 
+ WL[192] WL[193] WL[194] WL[195] WLPY[3] WLPYB[3] NET64[0] NET63[0] NET62[0] 
+ S1AHSF400W40_WLDV_2X1
XWLDV_2X1<49> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] NET68[4] 
+ NET68[5] NET68[6] NET68[7] NET67[8] NET67[9] NET67[10] NET67[11] NET67[12] 
+ NET67[13] NET67[14] NET67[15] NET66[8] NET66[9] NET66[10] NET66[11] 
+ NET66[12] NET66[13] NET66[14] NET66[15] PD_BUF PD_CVDDBUF NET65[1] VDDHD 
+ VDDI VSSI WL[196] WL[197] WL[198] WL[199] WLPY[3] WLPYB[3] NET64[1] NET63[1] 
+ NET62[1] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<50> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[1] NET68[8] 
+ NET68[9] NET68[10] NET68[11] NET67[16] NET67[17] NET67[18] NET67[19] 
+ NET67[20] NET67[21] NET67[22] NET67[23] NET66[16] NET66[17] NET66[18] 
+ NET66[19] NET66[20] NET66[21] NET66[22] NET66[23] PD_BUF PD_CVDDBUF NET65[2] 
+ VDDHD VDDI VSSI WL[200] WL[201] WL[202] WL[203] WLPY[3] WLPYB[3] NET64[2] 
+ NET63[2] NET62[2] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<51> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[1] NET68[12] 
+ NET68[13] NET68[14] NET68[15] NET67[24] NET67[25] NET67[26] NET67[27] 
+ NET67[28] NET67[29] NET67[30] NET67[31] NET66[24] NET66[25] NET66[26] 
+ NET66[27] NET66[28] NET66[29] NET66[30] NET66[31] PD_BUF PD_CVDDBUF NET65[3] 
+ VDDHD VDDI VSSI WL[204] WL[205] WL[206] WL[207] WLPY[3] WLPYB[3] NET64[3] 
+ NET63[3] NET62[3] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<52> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[2] NET68[16] 
+ NET68[17] NET68[18] NET68[19] NET67[32] NET67[33] NET67[34] NET67[35] 
+ NET67[36] NET67[37] NET67[38] NET67[39] NET66[32] NET66[33] NET66[34] 
+ NET66[35] NET66[36] NET66[37] NET66[38] NET66[39] PD_BUF PD_CVDDBUF NET65[4] 
+ VDDHD VDDI VSSI WL[208] WL[209] WL[210] WL[211] WLPY[3] WLPYB[3] NET64[4] 
+ NET63[4] NET62[4] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<53> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[2] NET68[20] 
+ NET68[21] NET68[22] NET68[23] NET67[40] NET67[41] NET67[42] NET67[43] 
+ NET67[44] NET67[45] NET67[46] NET67[47] NET66[40] NET66[41] NET66[42] 
+ NET66[43] NET66[44] NET66[45] NET66[46] NET66[47] PD_BUF PD_CVDDBUF NET65[5] 
+ VDDHD VDDI VSSI WL[212] WL[213] WL[214] WL[215] WLPY[3] WLPYB[3] NET64[5] 
+ NET63[5] NET62[5] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<54> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[3] NET68[24] 
+ NET68[25] NET68[26] NET68[27] NET67[48] NET67[49] NET67[50] NET67[51] 
+ NET67[52] NET67[53] NET67[54] NET67[55] NET66[48] NET66[49] NET66[50] 
+ NET66[51] NET66[52] NET66[53] NET66[54] NET66[55] PD_BUF PD_CVDDBUF NET65[6] 
+ VDDHD VDDI VSSI WL[216] WL[217] WL[218] WL[219] WLPY[3] WLPYB[3] NET64[6] 
+ NET63[6] NET62[6] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<55> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[3] NET68[28] 
+ NET68[29] NET68[30] NET68[31] NET67[56] NET67[57] NET67[58] NET67[59] 
+ NET67[60] NET67[61] NET67[62] NET67[63] NET66[56] NET66[57] NET66[58] 
+ NET66[59] NET66[60] NET66[61] NET66[62] NET66[63] PD_BUF PD_CVDDBUF NET65[7] 
+ VDDHD VDDI VSSI WL[220] WL[221] WL[222] WL[223] WLPY[3] WLPYB[3] NET64[7] 
+ NET63[7] NET62[7] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<56> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[4] NET68[32] 
+ NET68[33] NET68[34] NET68[35] NET67[64] NET67[65] NET67[66] NET67[67] 
+ NET67[68] NET67[69] NET67[70] NET67[71] NET66[64] NET66[65] NET66[66] 
+ NET66[67] NET66[68] NET66[69] NET66[70] NET66[71] PD_BUF PD_CVDDBUF NET65[8] 
+ VDDHD VDDI VSSI WL[224] WL[225] WL[226] WL[227] WLPY[3] WLPYB[3] NET64[8] 
+ NET63[8] NET62[8] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<57> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[4] NET68[36] 
+ NET68[37] NET68[38] NET68[39] NET67[72] NET67[73] NET67[74] NET67[75] 
+ NET67[76] NET67[77] NET67[78] NET67[79] NET66[72] NET66[73] NET66[74] 
+ NET66[75] NET66[76] NET66[77] NET66[78] NET66[79] PD_BUF PD_CVDDBUF NET65[9] 
+ VDDHD VDDI VSSI WL[228] WL[229] WL[230] WL[231] WLPY[3] WLPYB[3] NET64[9] 
+ NET63[9] NET62[9] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<58> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[5] NET68[40] 
+ NET68[41] NET68[42] NET68[43] NET67[80] NET67[81] NET67[82] NET67[83] 
+ NET67[84] NET67[85] NET67[86] NET67[87] NET66[80] NET66[81] NET66[82] 
+ NET66[83] NET66[84] NET66[85] NET66[86] NET66[87] PD_BUF PD_CVDDBUF 
+ NET65[10] VDDHD VDDI VSSI WL[232] WL[233] WL[234] WL[235] WLPY[3] WLPYB[3] 
+ NET64[10] NET63[10] NET62[10] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<59> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[5] NET68[44] 
+ NET68[45] NET68[46] NET68[47] NET67[88] NET67[89] NET67[90] NET67[91] 
+ NET67[92] NET67[93] NET67[94] NET67[95] NET66[88] NET66[89] NET66[90] 
+ NET66[91] NET66[92] NET66[93] NET66[94] NET66[95] PD_BUF PD_CVDDBUF 
+ NET65[11] VDDHD VDDI VSSI WL[236] WL[237] WL[238] WL[239] WLPY[3] WLPYB[3] 
+ NET64[11] NET63[11] NET62[11] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<60> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[6] NET68[48] 
+ NET68[49] NET68[50] NET68[51] NET67[96] NET67[97] NET67[98] NET67[99] 
+ NET67[100] NET67[101] NET67[102] NET67[103] NET66[96] NET66[97] NET66[98] 
+ NET66[99] NET66[100] NET66[101] NET66[102] NET66[103] PD_BUF PD_CVDDBUF 
+ NET65[12] VDDHD VDDI VSSI WL[240] WL[241] WL[242] WL[243] WLPY[3] WLPYB[3] 
+ NET64[12] NET63[12] NET62[12] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<61> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[6] NET68[52] 
+ NET68[53] NET68[54] NET68[55] NET67[104] NET67[105] NET67[106] NET67[107] 
+ NET67[108] NET67[109] NET67[110] NET67[111] NET66[104] NET66[105] NET66[106] 
+ NET66[107] NET66[108] NET66[109] NET66[110] NET66[111] PD_BUF PD_CVDDBUF 
+ NET65[13] VDDHD VDDI VSSI WL[244] WL[245] WL[246] WL[247] WLPY[3] WLPYB[3] 
+ NET64[13] NET63[13] NET62[13] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<62> DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X1[7] NET68[56] 
+ NET68[57] NET68[58] NET68[59] NET67[112] NET67[113] NET67[114] NET67[115] 
+ NET67[116] NET67[117] NET67[118] NET67[119] NET66[112] NET66[113] NET66[114] 
+ NET66[115] NET66[116] NET66[117] NET66[118] NET66[119] PD_BUF PD_CVDDBUF 
+ NET65[14] VDDHD VDDI VSSI WL[248] WL[249] WL[250] WL[251] WLPY[3] WLPYB[3] 
+ NET64[14] NET63[14] NET62[14] S1AHSF400W40_WLDV_2X1
XWLDV_2X1<63> DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[7] NET68[60] 
+ NET68[61] NET68[62] NET68[63] NET67[120] NET67[121] NET67[122] NET67[123] 
+ NET67[124] NET67[125] NET67[126] NET67[127] NET66[120] NET66[121] NET66[122] 
+ NET66[123] NET66[124] NET66[125] NET66[126] NET66[127] PD_BUF PD_CVDDBUF 
+ NET65[15] VDDHD VDDI VSSI WL[252] WL[253] WL[254] WL[255] WLPY[3] WLPYB[3] 
+ NET64[15] NET63[15] NET62[15] S1AHSF400W40_WLDV_2X1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_LCNT2_SEG6_S256
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_LCNT2_SEG6_S256 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] 
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] PD_BUF RW_RE VDDHD VDDI VSSI WLP_SAE WLP_SAE_TK YL[0]
*.PININFO DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B 
*.PININFO DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B 
*.PININFO DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B 
*.PININFO DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B DEC_X2[3]:B 
*.PININFO DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B DEC_X3[4]:B 
*.PININFO DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B DEC_Y[1]:B DEC_Y[2]:B 
*.PININFO DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B DEC_Y[7]:B PD_BUF:B 
*.PININFO RW_RE:B VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XI4 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] PD_BUF NET045 VDDHD VDDI VSSI NET37[0] NET37[1] NET37[2] 
+ NET37[3] NET37[4] NET37[5] NET37[6] NET37[7] NET37[8] NET37[9] NET37[10] 
+ NET37[11] NET37[12] NET37[13] NET37[14] NET37[15] NET37[16] NET37[17] 
+ NET37[18] NET37[19] NET37[20] NET37[21] NET37[22] NET37[23] NET37[24] 
+ NET37[25] NET37[26] NET37[27] NET37[28] NET37[29] NET37[30] NET37[31] 
+ NET37[32] NET37[33] NET37[34] NET37[35] NET37[36] NET37[37] NET37[38] 
+ NET37[39] NET37[40] NET37[41] NET37[42] NET37[43] NET37[44] NET37[45] 
+ NET37[46] NET37[47] NET37[48] NET37[49] NET37[50] NET37[51] NET37[52] 
+ NET37[53] NET37[54] NET37[55] NET37[56] NET37[57] NET37[58] NET37[59] 
+ NET37[60] NET37[61] NET37[62] NET37[63] NET37[64] NET37[65] NET37[66] 
+ NET37[67] NET37[68] NET37[69] NET37[70] NET37[71] NET37[72] NET37[73] 
+ NET37[74] NET37[75] NET37[76] NET37[77] NET37[78] NET37[79] NET37[80] 
+ NET37[81] NET37[82] NET37[83] NET37[84] NET37[85] NET37[86] NET37[87] 
+ NET37[88] NET37[89] NET37[90] NET37[91] NET37[92] NET37[93] NET37[94] 
+ NET37[95] NET37[96] NET37[97] NET37[98] NET37[99] NET37[100] NET37[101] 
+ NET37[102] NET37[103] NET37[104] NET37[105] NET37[106] NET37[107] NET37[108] 
+ NET37[109] NET37[110] NET37[111] NET37[112] NET37[113] NET37[114] NET37[115] 
+ NET37[116] NET37[117] NET37[118] NET37[119] NET37[120] NET37[121] NET37[122] 
+ NET37[123] NET37[124] NET37[125] NET37[126] NET37[127] NET37[128] NET37[129] 
+ NET37[130] NET37[131] NET37[132] NET37[133] NET37[134] NET37[135] NET37[136] 
+ NET37[137] NET37[138] NET37[139] NET37[140] NET37[141] NET37[142] NET37[143] 
+ NET37[144] NET37[145] NET37[146] NET37[147] NET37[148] NET37[149] NET37[150] 
+ NET37[151] NET37[152] NET37[153] NET37[154] NET37[155] NET37[156] NET37[157] 
+ NET37[158] NET37[159] NET37[160] NET37[161] NET37[162] NET37[163] NET37[164] 
+ NET37[165] NET37[166] NET37[167] NET37[168] NET37[169] NET37[170] NET37[171] 
+ NET37[172] NET37[173] NET37[174] NET37[175] NET37[176] NET37[177] NET37[178] 
+ NET37[179] NET37[180] NET37[181] NET37[182] NET37[183] NET37[184] NET37[185] 
+ NET37[186] NET37[187] NET37[188] NET37[189] NET37[190] NET37[191] NET37[192] 
+ NET37[193] NET37[194] NET37[195] NET37[196] NET37[197] NET37[198] NET37[199] 
+ NET37[200] NET37[201] NET37[202] NET37[203] NET37[204] NET37[205] NET37[206] 
+ NET37[207] NET37[208] NET37[209] NET37[210] NET37[211] NET37[212] NET37[213] 
+ NET37[214] NET37[215] NET37[216] NET37[217] NET37[218] NET37[219] NET37[220] 
+ NET37[221] NET37[222] NET37[223] NET37[224] NET37[225] NET37[226] NET37[227] 
+ NET37[228] NET37[229] NET37[230] NET37[231] NET37[232] NET37[233] NET37[234] 
+ NET37[235] NET37[236] NET37[237] NET37[238] NET37[239] NET37[240] NET37[241] 
+ NET37[242] NET37[243] NET37[244] NET37[245] NET37[246] NET37[247] NET37[248] 
+ NET37[249] NET37[250] NET37[251] NET37[252] NET37[253] NET37[254] NET37[255] 
+ WLPY_0UP[0] WLPY_0UP[1] WLPY_0UP[2] WLPY_0UP[3] WLPYB_0UP[0] WLPYB_0UP[1] 
+ WLPYB_0UP[2] WLPYB_0UP[3] S1AHSF400W40_WLDV_256X1
XI3 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] PD_BUF NET055 VDDHD VDDI VSSI NET47[0] NET47[1] NET47[2] 
+ NET47[3] NET47[4] NET47[5] NET47[6] NET47[7] NET47[8] NET47[9] NET47[10] 
+ NET47[11] NET47[12] NET47[13] NET47[14] NET47[15] NET47[16] NET47[17] 
+ NET47[18] NET47[19] NET47[20] NET47[21] NET47[22] NET47[23] NET47[24] 
+ NET47[25] NET47[26] NET47[27] NET47[28] NET47[29] NET47[30] NET47[31] 
+ NET47[32] NET47[33] NET47[34] NET47[35] NET47[36] NET47[37] NET47[38] 
+ NET47[39] NET47[40] NET47[41] NET47[42] NET47[43] NET47[44] NET47[45] 
+ NET47[46] NET47[47] NET47[48] NET47[49] NET47[50] NET47[51] NET47[52] 
+ NET47[53] NET47[54] NET47[55] NET47[56] NET47[57] NET47[58] NET47[59] 
+ NET47[60] NET47[61] NET47[62] NET47[63] NET47[64] NET47[65] NET47[66] 
+ NET47[67] NET47[68] NET47[69] NET47[70] NET47[71] NET47[72] NET47[73] 
+ NET47[74] NET47[75] NET47[76] NET47[77] NET47[78] NET47[79] NET47[80] 
+ NET47[81] NET47[82] NET47[83] NET47[84] NET47[85] NET47[86] NET47[87] 
+ NET47[88] NET47[89] NET47[90] NET47[91] NET47[92] NET47[93] NET47[94] 
+ NET47[95] NET47[96] NET47[97] NET47[98] NET47[99] NET47[100] NET47[101] 
+ NET47[102] NET47[103] NET47[104] NET47[105] NET47[106] NET47[107] NET47[108] 
+ NET47[109] NET47[110] NET47[111] NET47[112] NET47[113] NET47[114] NET47[115] 
+ NET47[116] NET47[117] NET47[118] NET47[119] NET47[120] NET47[121] NET47[122] 
+ NET47[123] NET47[124] NET47[125] NET47[126] NET47[127] NET47[128] NET47[129] 
+ NET47[130] NET47[131] NET47[132] NET47[133] NET47[134] NET47[135] NET47[136] 
+ NET47[137] NET47[138] NET47[139] NET47[140] NET47[141] NET47[142] NET47[143] 
+ NET47[144] NET47[145] NET47[146] NET47[147] NET47[148] NET47[149] NET47[150] 
+ NET47[151] NET47[152] NET47[153] NET47[154] NET47[155] NET47[156] NET47[157] 
+ NET47[158] NET47[159] NET47[160] NET47[161] NET47[162] NET47[163] NET47[164] 
+ NET47[165] NET47[166] NET47[167] NET47[168] NET47[169] NET47[170] NET47[171] 
+ NET47[172] NET47[173] NET47[174] NET47[175] NET47[176] NET47[177] NET47[178] 
+ NET47[179] NET47[180] NET47[181] NET47[182] NET47[183] NET47[184] NET47[185] 
+ NET47[186] NET47[187] NET47[188] NET47[189] NET47[190] NET47[191] NET47[192] 
+ NET47[193] NET47[194] NET47[195] NET47[196] NET47[197] NET47[198] NET47[199] 
+ NET47[200] NET47[201] NET47[202] NET47[203] NET47[204] NET47[205] NET47[206] 
+ NET47[207] NET47[208] NET47[209] NET47[210] NET47[211] NET47[212] NET47[213] 
+ NET47[214] NET47[215] NET47[216] NET47[217] NET47[218] NET47[219] NET47[220] 
+ NET47[221] NET47[222] NET47[223] NET47[224] NET47[225] NET47[226] NET47[227] 
+ NET47[228] NET47[229] NET47[230] NET47[231] NET47[232] NET47[233] NET47[234] 
+ NET47[235] NET47[236] NET47[237] NET47[238] NET47[239] NET47[240] NET47[241] 
+ NET47[242] NET47[243] NET47[244] NET47[245] NET47[246] NET47[247] NET47[248] 
+ NET47[249] NET47[250] NET47[251] NET47[252] NET47[253] NET47[254] NET47[255] 
+ WLPY_3DN[0] WLPY_3DN[1] WLPY_3DN[2] WLPY_3DN[3] WLPYB_3DN[0] WLPYB_3DN[1] 
+ WLPYB_3DN[2] WLPYB_3DN[3] S1AHSF400W40_WLDV_256X1
XI1 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] PD_BUF NET065 VDDHD VDDI VSSI NET57[0] NET57[1] NET57[2] 
+ NET57[3] NET57[4] NET57[5] NET57[6] NET57[7] NET57[8] NET57[9] NET57[10] 
+ NET57[11] NET57[12] NET57[13] NET57[14] NET57[15] NET57[16] NET57[17] 
+ NET57[18] NET57[19] NET57[20] NET57[21] NET57[22] NET57[23] NET57[24] 
+ NET57[25] NET57[26] NET57[27] NET57[28] NET57[29] NET57[30] NET57[31] 
+ NET57[32] NET57[33] NET57[34] NET57[35] NET57[36] NET57[37] NET57[38] 
+ NET57[39] NET57[40] NET57[41] NET57[42] NET57[43] NET57[44] NET57[45] 
+ NET57[46] NET57[47] NET57[48] NET57[49] NET57[50] NET57[51] NET57[52] 
+ NET57[53] NET57[54] NET57[55] NET57[56] NET57[57] NET57[58] NET57[59] 
+ NET57[60] NET57[61] NET57[62] NET57[63] NET57[64] NET57[65] NET57[66] 
+ NET57[67] NET57[68] NET57[69] NET57[70] NET57[71] NET57[72] NET57[73] 
+ NET57[74] NET57[75] NET57[76] NET57[77] NET57[78] NET57[79] NET57[80] 
+ NET57[81] NET57[82] NET57[83] NET57[84] NET57[85] NET57[86] NET57[87] 
+ NET57[88] NET57[89] NET57[90] NET57[91] NET57[92] NET57[93] NET57[94] 
+ NET57[95] NET57[96] NET57[97] NET57[98] NET57[99] NET57[100] NET57[101] 
+ NET57[102] NET57[103] NET57[104] NET57[105] NET57[106] NET57[107] NET57[108] 
+ NET57[109] NET57[110] NET57[111] NET57[112] NET57[113] NET57[114] NET57[115] 
+ NET57[116] NET57[117] NET57[118] NET57[119] NET57[120] NET57[121] NET57[122] 
+ NET57[123] NET57[124] NET57[125] NET57[126] NET57[127] NET57[128] NET57[129] 
+ NET57[130] NET57[131] NET57[132] NET57[133] NET57[134] NET57[135] NET57[136] 
+ NET57[137] NET57[138] NET57[139] NET57[140] NET57[141] NET57[142] NET57[143] 
+ NET57[144] NET57[145] NET57[146] NET57[147] NET57[148] NET57[149] NET57[150] 
+ NET57[151] NET57[152] NET57[153] NET57[154] NET57[155] NET57[156] NET57[157] 
+ NET57[158] NET57[159] NET57[160] NET57[161] NET57[162] NET57[163] NET57[164] 
+ NET57[165] NET57[166] NET57[167] NET57[168] NET57[169] NET57[170] NET57[171] 
+ NET57[172] NET57[173] NET57[174] NET57[175] NET57[176] NET57[177] NET57[178] 
+ NET57[179] NET57[180] NET57[181] NET57[182] NET57[183] NET57[184] NET57[185] 
+ NET57[186] NET57[187] NET57[188] NET57[189] NET57[190] NET57[191] NET57[192] 
+ NET57[193] NET57[194] NET57[195] NET57[196] NET57[197] NET57[198] NET57[199] 
+ NET57[200] NET57[201] NET57[202] NET57[203] NET57[204] NET57[205] NET57[206] 
+ NET57[207] NET57[208] NET57[209] NET57[210] NET57[211] NET57[212] NET57[213] 
+ NET57[214] NET57[215] NET57[216] NET57[217] NET57[218] NET57[219] NET57[220] 
+ NET57[221] NET57[222] NET57[223] NET57[224] NET57[225] NET57[226] NET57[227] 
+ NET57[228] NET57[229] NET57[230] NET57[231] NET57[232] NET57[233] NET57[234] 
+ NET57[235] NET57[236] NET57[237] NET57[238] NET57[239] NET57[240] NET57[241] 
+ NET57[242] NET57[243] NET57[244] NET57[245] NET57[246] NET57[247] NET57[248] 
+ NET57[249] NET57[250] NET57[251] NET57[252] NET57[253] NET57[254] NET57[255] 
+ WLPY_1DN[0] WLPY_1DN[1] WLPY_1DN[2] WLPY_1DN[3] WLPYB_1DN[0] WLPYB_1DN[1] 
+ WLPYB_1DN[2] WLPYB_1DN[3] S1AHSF400W40_WLDV_256X1
XI0 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] PD_BUF NET075 VDDHD VDDI VSSI NET67[0] NET67[1] NET67[2] 
+ NET67[3] NET67[4] NET67[5] NET67[6] NET67[7] NET67[8] NET67[9] NET67[10] 
+ NET67[11] NET67[12] NET67[13] NET67[14] NET67[15] NET67[16] NET67[17] 
+ NET67[18] NET67[19] NET67[20] NET67[21] NET67[22] NET67[23] NET67[24] 
+ NET67[25] NET67[26] NET67[27] NET67[28] NET67[29] NET67[30] NET67[31] 
+ NET67[32] NET67[33] NET67[34] NET67[35] NET67[36] NET67[37] NET67[38] 
+ NET67[39] NET67[40] NET67[41] NET67[42] NET67[43] NET67[44] NET67[45] 
+ NET67[46] NET67[47] NET67[48] NET67[49] NET67[50] NET67[51] NET67[52] 
+ NET67[53] NET67[54] NET67[55] NET67[56] NET67[57] NET67[58] NET67[59] 
+ NET67[60] NET67[61] NET67[62] NET67[63] NET67[64] NET67[65] NET67[66] 
+ NET67[67] NET67[68] NET67[69] NET67[70] NET67[71] NET67[72] NET67[73] 
+ NET67[74] NET67[75] NET67[76] NET67[77] NET67[78] NET67[79] NET67[80] 
+ NET67[81] NET67[82] NET67[83] NET67[84] NET67[85] NET67[86] NET67[87] 
+ NET67[88] NET67[89] NET67[90] NET67[91] NET67[92] NET67[93] NET67[94] 
+ NET67[95] NET67[96] NET67[97] NET67[98] NET67[99] NET67[100] NET67[101] 
+ NET67[102] NET67[103] NET67[104] NET67[105] NET67[106] NET67[107] NET67[108] 
+ NET67[109] NET67[110] NET67[111] NET67[112] NET67[113] NET67[114] NET67[115] 
+ NET67[116] NET67[117] NET67[118] NET67[119] NET67[120] NET67[121] NET67[122] 
+ NET67[123] NET67[124] NET67[125] NET67[126] NET67[127] NET67[128] NET67[129] 
+ NET67[130] NET67[131] NET67[132] NET67[133] NET67[134] NET67[135] NET67[136] 
+ NET67[137] NET67[138] NET67[139] NET67[140] NET67[141] NET67[142] NET67[143] 
+ NET67[144] NET67[145] NET67[146] NET67[147] NET67[148] NET67[149] NET67[150] 
+ NET67[151] NET67[152] NET67[153] NET67[154] NET67[155] NET67[156] NET67[157] 
+ NET67[158] NET67[159] NET67[160] NET67[161] NET67[162] NET67[163] NET67[164] 
+ NET67[165] NET67[166] NET67[167] NET67[168] NET67[169] NET67[170] NET67[171] 
+ NET67[172] NET67[173] NET67[174] NET67[175] NET67[176] NET67[177] NET67[178] 
+ NET67[179] NET67[180] NET67[181] NET67[182] NET67[183] NET67[184] NET67[185] 
+ NET67[186] NET67[187] NET67[188] NET67[189] NET67[190] NET67[191] NET67[192] 
+ NET67[193] NET67[194] NET67[195] NET67[196] NET67[197] NET67[198] NET67[199] 
+ NET67[200] NET67[201] NET67[202] NET67[203] NET67[204] NET67[205] NET67[206] 
+ NET67[207] NET67[208] NET67[209] NET67[210] NET67[211] NET67[212] NET67[213] 
+ NET67[214] NET67[215] NET67[216] NET67[217] NET67[218] NET67[219] NET67[220] 
+ NET67[221] NET67[222] NET67[223] NET67[224] NET67[225] NET67[226] NET67[227] 
+ NET67[228] NET67[229] NET67[230] NET67[231] NET67[232] NET67[233] NET67[234] 
+ NET67[235] NET67[236] NET67[237] NET67[238] NET67[239] NET67[240] NET67[241] 
+ NET67[242] NET67[243] NET67[244] NET67[245] NET67[246] NET67[247] NET67[248] 
+ NET67[249] NET67[250] NET67[251] NET67[252] NET67[253] NET67[254] NET67[255] 
+ WLPY_1UP[0] WLPY_1UP[1] WLPY_1UP[2] WLPY_1UP[3] WLPYB_1UP[0] WLPYB_1UP[1] 
+ WLPYB_1UP[2] WLPYB_1UP[3] S1AHSF400W40_WLDV_256X1
XWLDV_256X1_U DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] PD_BUF NET085 VDDHD VDDI VSSI NET77[0] 
+ NET77[1] NET77[2] NET77[3] NET77[4] NET77[5] NET77[6] NET77[7] NET77[8] 
+ NET77[9] NET77[10] NET77[11] NET77[12] NET77[13] NET77[14] NET77[15] 
+ NET77[16] NET77[17] NET77[18] NET77[19] NET77[20] NET77[21] NET77[22] 
+ NET77[23] NET77[24] NET77[25] NET77[26] NET77[27] NET77[28] NET77[29] 
+ NET77[30] NET77[31] NET77[32] NET77[33] NET77[34] NET77[35] NET77[36] 
+ NET77[37] NET77[38] NET77[39] NET77[40] NET77[41] NET77[42] NET77[43] 
+ NET77[44] NET77[45] NET77[46] NET77[47] NET77[48] NET77[49] NET77[50] 
+ NET77[51] NET77[52] NET77[53] NET77[54] NET77[55] NET77[56] NET77[57] 
+ NET77[58] NET77[59] NET77[60] NET77[61] NET77[62] NET77[63] NET77[64] 
+ NET77[65] NET77[66] NET77[67] NET77[68] NET77[69] NET77[70] NET77[71] 
+ NET77[72] NET77[73] NET77[74] NET77[75] NET77[76] NET77[77] NET77[78] 
+ NET77[79] NET77[80] NET77[81] NET77[82] NET77[83] NET77[84] NET77[85] 
+ NET77[86] NET77[87] NET77[88] NET77[89] NET77[90] NET77[91] NET77[92] 
+ NET77[93] NET77[94] NET77[95] NET77[96] NET77[97] NET77[98] NET77[99] 
+ NET77[100] NET77[101] NET77[102] NET77[103] NET77[104] NET77[105] NET77[106] 
+ NET77[107] NET77[108] NET77[109] NET77[110] NET77[111] NET77[112] NET77[113] 
+ NET77[114] NET77[115] NET77[116] NET77[117] NET77[118] NET77[119] NET77[120] 
+ NET77[121] NET77[122] NET77[123] NET77[124] NET77[125] NET77[126] NET77[127] 
+ NET77[128] NET77[129] NET77[130] NET77[131] NET77[132] NET77[133] NET77[134] 
+ NET77[135] NET77[136] NET77[137] NET77[138] NET77[139] NET77[140] NET77[141] 
+ NET77[142] NET77[143] NET77[144] NET77[145] NET77[146] NET77[147] NET77[148] 
+ NET77[149] NET77[150] NET77[151] NET77[152] NET77[153] NET77[154] NET77[155] 
+ NET77[156] NET77[157] NET77[158] NET77[159] NET77[160] NET77[161] NET77[162] 
+ NET77[163] NET77[164] NET77[165] NET77[166] NET77[167] NET77[168] NET77[169] 
+ NET77[170] NET77[171] NET77[172] NET77[173] NET77[174] NET77[175] NET77[176] 
+ NET77[177] NET77[178] NET77[179] NET77[180] NET77[181] NET77[182] NET77[183] 
+ NET77[184] NET77[185] NET77[186] NET77[187] NET77[188] NET77[189] NET77[190] 
+ NET77[191] NET77[192] NET77[193] NET77[194] NET77[195] NET77[196] NET77[197] 
+ NET77[198] NET77[199] NET77[200] NET77[201] NET77[202] NET77[203] NET77[204] 
+ NET77[205] NET77[206] NET77[207] NET77[208] NET77[209] NET77[210] NET77[211] 
+ NET77[212] NET77[213] NET77[214] NET77[215] NET77[216] NET77[217] NET77[218] 
+ NET77[219] NET77[220] NET77[221] NET77[222] NET77[223] NET77[224] NET77[225] 
+ NET77[226] NET77[227] NET77[228] NET77[229] NET77[230] NET77[231] NET77[232] 
+ NET77[233] NET77[234] NET77[235] NET77[236] NET77[237] NET77[238] NET77[239] 
+ NET77[240] NET77[241] NET77[242] NET77[243] NET77[244] NET77[245] NET77[246] 
+ NET77[247] NET77[248] NET77[249] NET77[250] NET77[251] NET77[252] NET77[253] 
+ NET77[254] NET77[255] WLPY_2UP[0] WLPY_2UP[1] WLPY_2UP[2] WLPY_2UP[3] 
+ WLPYB_2UP[0] WLPYB_2UP[1] WLPYB_2UP[2] WLPYB_2UP[3] S1AHSF400W40_WLDV_256X1
XWLDV_256X1_D DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] 
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] PD_BUF NET095 VDDHD VDDI VSSI NET87[0] 
+ NET87[1] NET87[2] NET87[3] NET87[4] NET87[5] NET87[6] NET87[7] NET87[8] 
+ NET87[9] NET87[10] NET87[11] NET87[12] NET87[13] NET87[14] NET87[15] 
+ NET87[16] NET87[17] NET87[18] NET87[19] NET87[20] NET87[21] NET87[22] 
+ NET87[23] NET87[24] NET87[25] NET87[26] NET87[27] NET87[28] NET87[29] 
+ NET87[30] NET87[31] NET87[32] NET87[33] NET87[34] NET87[35] NET87[36] 
+ NET87[37] NET87[38] NET87[39] NET87[40] NET87[41] NET87[42] NET87[43] 
+ NET87[44] NET87[45] NET87[46] NET87[47] NET87[48] NET87[49] NET87[50] 
+ NET87[51] NET87[52] NET87[53] NET87[54] NET87[55] NET87[56] NET87[57] 
+ NET87[58] NET87[59] NET87[60] NET87[61] NET87[62] NET87[63] NET87[64] 
+ NET87[65] NET87[66] NET87[67] NET87[68] NET87[69] NET87[70] NET87[71] 
+ NET87[72] NET87[73] NET87[74] NET87[75] NET87[76] NET87[77] NET87[78] 
+ NET87[79] NET87[80] NET87[81] NET87[82] NET87[83] NET87[84] NET87[85] 
+ NET87[86] NET87[87] NET87[88] NET87[89] NET87[90] NET87[91] NET87[92] 
+ NET87[93] NET87[94] NET87[95] NET87[96] NET87[97] NET87[98] NET87[99] 
+ NET87[100] NET87[101] NET87[102] NET87[103] NET87[104] NET87[105] NET87[106] 
+ NET87[107] NET87[108] NET87[109] NET87[110] NET87[111] NET87[112] NET87[113] 
+ NET87[114] NET87[115] NET87[116] NET87[117] NET87[118] NET87[119] NET87[120] 
+ NET87[121] NET87[122] NET87[123] NET87[124] NET87[125] NET87[126] NET87[127] 
+ NET87[128] NET87[129] NET87[130] NET87[131] NET87[132] NET87[133] NET87[134] 
+ NET87[135] NET87[136] NET87[137] NET87[138] NET87[139] NET87[140] NET87[141] 
+ NET87[142] NET87[143] NET87[144] NET87[145] NET87[146] NET87[147] NET87[148] 
+ NET87[149] NET87[150] NET87[151] NET87[152] NET87[153] NET87[154] NET87[155] 
+ NET87[156] NET87[157] NET87[158] NET87[159] NET87[160] NET87[161] NET87[162] 
+ NET87[163] NET87[164] NET87[165] NET87[166] NET87[167] NET87[168] NET87[169] 
+ NET87[170] NET87[171] NET87[172] NET87[173] NET87[174] NET87[175] NET87[176] 
+ NET87[177] NET87[178] NET87[179] NET87[180] NET87[181] NET87[182] NET87[183] 
+ NET87[184] NET87[185] NET87[186] NET87[187] NET87[188] NET87[189] NET87[190] 
+ NET87[191] NET87[192] NET87[193] NET87[194] NET87[195] NET87[196] NET87[197] 
+ NET87[198] NET87[199] NET87[200] NET87[201] NET87[202] NET87[203] NET87[204] 
+ NET87[205] NET87[206] NET87[207] NET87[208] NET87[209] NET87[210] NET87[211] 
+ NET87[212] NET87[213] NET87[214] NET87[215] NET87[216] NET87[217] NET87[218] 
+ NET87[219] NET87[220] NET87[221] NET87[222] NET87[223] NET87[224] NET87[225] 
+ NET87[226] NET87[227] NET87[228] NET87[229] NET87[230] NET87[231] NET87[232] 
+ NET87[233] NET87[234] NET87[235] NET87[236] NET87[237] NET87[238] NET87[239] 
+ NET87[240] NET87[241] NET87[242] NET87[243] NET87[244] NET87[245] NET87[246] 
+ NET87[247] NET87[248] NET87[249] NET87[250] NET87[251] NET87[252] NET87[253] 
+ NET87[254] NET87[255] WLPY_2DN[0] WLPY_2DN[1] WLPY_2DN[2] WLPY_2DN[3] 
+ WLPYB_2DN[0] WLPYB_2DN[1] WLPYB_2DN[2] WLPYB_2DN[3] S1AHSF400W40_WLDV_256X1
XXDRV_STRP_1D<0> VDDHD VDDI VSSI WLPY_1DN[0] WLPYB_1DN[0] S1AHSF400W40_XDRV_STRAP
XXDRV_STRP_1D<1> VDDHD VDDI VSSI WLPY_1DN[1] WLPYB_1DN[1] S1AHSF400W40_XDRV_STRAP
XXDRV_STRP_1D<2> VDDHD VDDI VSSI WLPY_1DN[2] WLPYB_1DN[2] S1AHSF400W40_XDRV_STRAP
XXDRV_STRP_1D<3> VDDHD VDDI VSSI WLPY_1DN[3] WLPYB_1DN[3] S1AHSF400W40_XDRV_STRAP
XI7<0> VDDHD VDDI VSSI WLPY_2UP[0] WLPYB_2UP[0] S1AHSF400W40_XDRV_STRAP
XI7<1> VDDHD VDDI VSSI WLPY_2UP[1] WLPYB_2UP[1] S1AHSF400W40_XDRV_STRAP
XI7<2> VDDHD VDDI VSSI WLPY_2UP[2] WLPYB_2UP[2] S1AHSF400W40_XDRV_STRAP
XI7<3> VDDHD VDDI VSSI WLPY_2UP[3] WLPYB_2UP[3] S1AHSF400W40_XDRV_STRAP
XI6<0> VDDHD VDDI VSSI WLPY_2DN[0] WLPYB_2DN[0] S1AHSF400W40_XDRV_STRAP
XI6<1> VDDHD VDDI VSSI WLPY_2DN[1] WLPYB_2DN[1] S1AHSF400W40_XDRV_STRAP
XI6<2> VDDHD VDDI VSSI WLPY_2DN[2] WLPYB_2DN[2] S1AHSF400W40_XDRV_STRAP
XI6<3> VDDHD VDDI VSSI WLPY_2DN[3] WLPYB_2DN[3] S1AHSF400W40_XDRV_STRAP
XXDRV_STRAP_1U<0> VDDHD VDDI VSSI WLPY_1UP[0] WLPYB_1UP[0] S1AHSF400W40_XDRV_STRAP
XXDRV_STRAP_1U<1> VDDHD VDDI VSSI WLPY_1UP[1] WLPYB_1UP[1] S1AHSF400W40_XDRV_STRAP
XXDRV_STRAP_1U<2> VDDHD VDDI VSSI WLPY_1UP[2] WLPYB_1UP[2] S1AHSF400W40_XDRV_STRAP
XXDRV_STRAP_1U<3> VDDHD VDDI VSSI WLPY_1UP[3] WLPYB_1UP[3] S1AHSF400W40_XDRV_STRAP
XI2 NET108 NET106 NET0117[0] NET0117[1] NET0117[2] NET0117[3] NET0117[4] 
+ NET0117[5] NET0117[6] NET0117[7] NET0118[0] NET0118[1] NET0118[2] NET0118[3] 
+ NET0118[4] NET0118[5] NET0118[6] NET0118[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[2] DEC_X3[3] NET0116[0] NET0116[1] NET0116[2] NET0116[3] 
+ NET0116[4] NET0116[5] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] NET104[0] NET104[1] NET104[2] NET104[3] NET104[4] 
+ NET104[5] NET104[6] NET104[7] NET109[0] NET109[1] NET109[2] NET109[3] 
+ NET109[4] NET109[5] NET109[6] NET109[7] PD_BUF NET0103 NET110 RW_RE NET105 
+ VDDHD VDDI VSSI NET107 WLPY_1DN[0] WLPY_1DN[1] WLPY_1DN[2] WLPY_1DN[3] 
+ WLPY_1UP[0] WLPY_1UP[1] WLPY_1UP[2] WLPY_1UP[3] WLP_SAE NET0115 YL[0] 
+ NET95[0] NET95[1] S1AHSF400W40_LCTRL_S_M4
XLCTRL_S_M4 NET130 NET128 NET0142[0] NET0142[1] NET0142[2] NET0142[3] 
+ NET0142[4] NET0142[5] NET0142[6] NET0142[7] NET0143[0] NET0143[1] NET0143[2] 
+ NET0143[3] NET0143[4] NET0143[5] NET0143[6] NET0143[7] DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] DEC_X3[4] DEC_X3[5] NET0141[0] NET0141[1] NET0141[2] 
+ NET0141[3] NET0141[4] NET0141[5] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] 
+ DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] NET126[0] NET126[1] NET126[2] NET126[3] 
+ NET126[4] NET126[5] NET126[6] NET126[7] NET131[0] NET131[1] NET131[2] 
+ NET131[3] NET131[4] NET131[5] NET131[6] NET131[7] PD_BUF NET0125 NET132 
+ RW_RE NET127 VDDHD VDDI VSSI NET129 WLPY_2DN[0] WLPY_2DN[1] WLPY_2DN[2] 
+ WLPY_2DN[3] WLPY_2UP[0] WLPY_2UP[1] WLPY_2UP[2] WLPY_2UP[3] WLP_SAE NET011 
+ YL[0] NET117[0] NET117[1] S1AHSF400W40_LCTRL_S_M4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    BK_SEG_LD_SIM
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_BK_SEG_LD_SIM CVDDHD CVDDI DEC_X0_BT[0] DEC_X0_BT[1] DEC_X0_BT[2] 
+ DEC_X0_BT[3] DEC_X0_BT[4] DEC_X0_BT[5] DEC_X0_BT[6] DEC_X0_BT[7] 
+ DEC_X0_TP[0] DEC_X0_TP[1] DEC_X0_TP[2] DEC_X0_TP[3] DEC_X0_TP[4] 
+ DEC_X0_TP[5] DEC_X0_TP[6] DEC_X0_TP[7] DEC_X1_BT[0] DEC_X1_BT[1] 
+ DEC_X1_BT[2] DEC_X1_BT[3] DEC_X1_BT[4] DEC_X1_BT[5] DEC_X1_BT[6] 
+ DEC_X1_BT[7] DEC_X1_TP[0] DEC_X1_TP[1] DEC_X1_TP[2] DEC_X1_TP[3] 
+ DEC_X1_TP[4] DEC_X1_TP[5] DEC_X1_TP[6] DEC_X1_TP[7] DEC_X2_BT[0] 
+ DEC_X2_BT[1] DEC_X2_BT[2] DEC_X2_BT[3] DEC_X2_TP[0] DEC_X2_TP[1] 
+ DEC_X2_TP[2] DEC_X2_TP[3] DEC_X3_BT[0] DEC_X3_BT[1] DEC_X3_BT[2] 
+ DEC_X3_BT[3] DEC_X3_BT[4] DEC_X3_BT[5] DEC_X3_BT[6] DEC_X3_BT[7] 
+ DEC_X3_TP[0] DEC_X3_TP[1] DEC_X3_TP[2] DEC_X3_TP[3] DEC_X3_TP[4] 
+ DEC_X3_TP[5] DEC_X3_TP[6] DEC_X3_TP[7] DEC_Y_BT[0] DEC_Y_BT[1] DEC_Y_BT[2] 
+ DEC_Y_BT[3] DEC_Y_BT[4] DEC_Y_BT[5] DEC_Y_BT[6] DEC_Y_BT[7] DEC_Y_TP[0] 
+ DEC_Y_TP[1] DEC_Y_TP[2] DEC_Y_TP[3] DEC_Y_TP[4] DEC_Y_TP[5] DEC_Y_TP[6] 
+ DEC_Y_TP[7] PD_BUF_BT PD_BUF_TP PD_CVDDBUF_BT PD_CVDDBUF_TP RW_RE_BT 
+ RW_RE_TP VDDHD VDDI VSSI WLP_SAE_BT WLP_SAE_TK_BT WLP_SAE_TK_TP WLP_SAE_TP 
+ YL_BT[0] YL_TP[0]
*.PININFO DEC_X0_BT[0]:I DEC_X0_BT[1]:I DEC_X0_BT[2]:I DEC_X0_BT[3]:I 
*.PININFO DEC_X0_BT[4]:I DEC_X0_BT[5]:I DEC_X0_BT[6]:I DEC_X0_BT[7]:I 
*.PININFO DEC_X1_BT[0]:I DEC_X1_BT[1]:I DEC_X1_BT[2]:I DEC_X1_BT[3]:I 
*.PININFO DEC_X1_BT[4]:I DEC_X1_BT[5]:I DEC_X1_BT[6]:I DEC_X1_BT[7]:I 
*.PININFO PD_BUF_BT:I PD_CVDDBUF_BT:I RW_RE_TP:I DEC_X0_TP[0]:O DEC_X0_TP[1]:O 
*.PININFO DEC_X0_TP[2]:O DEC_X0_TP[3]:O DEC_X0_TP[4]:O DEC_X0_TP[5]:O 
*.PININFO DEC_X0_TP[6]:O DEC_X0_TP[7]:O DEC_X1_TP[0]:O DEC_X1_TP[1]:O 
*.PININFO DEC_X1_TP[2]:O DEC_X1_TP[3]:O DEC_X1_TP[4]:O DEC_X1_TP[5]:O 
*.PININFO DEC_X1_TP[6]:O DEC_X1_TP[7]:O PD_BUF_TP:O PD_CVDDBUF_TP:O CVDDHD:B 
*.PININFO CVDDI:B DEC_X2_BT[0]:B DEC_X2_BT[1]:B DEC_X2_BT[2]:B DEC_X2_BT[3]:B 
*.PININFO DEC_X2_TP[0]:B DEC_X2_TP[1]:B DEC_X2_TP[2]:B DEC_X2_TP[3]:B 
*.PININFO DEC_X3_BT[0]:B DEC_X3_BT[1]:B DEC_X3_BT[2]:B DEC_X3_BT[3]:B 
*.PININFO DEC_X3_BT[4]:B DEC_X3_BT[5]:B DEC_X3_BT[6]:B DEC_X3_BT[7]:B 
*.PININFO DEC_X3_TP[0]:B DEC_X3_TP[1]:B DEC_X3_TP[2]:B DEC_X3_TP[3]:B 
*.PININFO DEC_X3_TP[4]:B DEC_X3_TP[5]:B DEC_X3_TP[6]:B DEC_X3_TP[7]:B 
*.PININFO DEC_Y_BT[0]:B DEC_Y_BT[1]:B DEC_Y_BT[2]:B DEC_Y_BT[3]:B 
*.PININFO DEC_Y_BT[4]:B DEC_Y_BT[5]:B DEC_Y_BT[6]:B DEC_Y_BT[7]:B 
*.PININFO DEC_Y_TP[0]:B DEC_Y_TP[1]:B DEC_Y_TP[2]:B DEC_Y_TP[3]:B 
*.PININFO DEC_Y_TP[4]:B DEC_Y_TP[5]:B DEC_Y_TP[6]:B DEC_Y_TP[7]:B RW_RE_BT:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE_BT:B WLP_SAE_TK_BT:B WLP_SAE_TK_TP:B 
*.PININFO WLP_SAE_TP:B YL_BT[0]:B YL_TP[0]:B
XI25 NET039[0] NET039[1] NET039[2] NET039[3] NET039[4] NET039[5] NET039[6] 
+ NET039[7] NET036[0] NET036[1] NET036[2] NET036[3] NET036[4] NET036[5] 
+ NET036[6] NET036[7] NET034[0] NET034[1] NET034[2] NET034[3] NET033[0] 
+ NET033[1] NET033[2] NET033[3] NET033[4] NET033[5] NET033[6] NET033[7] 
+ NET032[0] NET032[1] NET032[2] NET032[3] NET032[4] NET032[5] NET032[6] 
+ NET032[7] NET031 NET035 NET037 NET040 NET041 NET030 NET029 NET03 
+ S1AHSF400W40_BK_LCNT2_SEG6_S64
XI24 NET39[0] NET39[1] NET39[2] NET39[3] NET39[4] NET39[5] NET39[6] NET39[7] 
+ NET36[0] NET36[1] NET36[2] NET36[3] NET36[4] NET36[5] NET36[6] NET36[7] 
+ NET34[0] NET34[1] NET34[2] NET34[3] NET33[0] NET33[1] NET33[2] NET33[3] 
+ NET33[4] NET33[5] NET33[6] NET33[7] NET32[0] NET32[1] NET32[2] NET32[3] 
+ NET32[4] NET32[5] NET32[6] NET32[7] NET31 NET35 NET37 NET40 NET41 NET30 
+ NET29 NET047 S1AHSF400W40_BK_LCNT2_SEG6_S256
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SIM_FULL
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SIM_FULL AWT BIST BWEBM_LL BWEBM_LR BWEB_LL BWEB_LR CEB CEBM CLK DM_LL 
+ DM_LR D_LL D_LR FAD1[0] FAD1[1] FAD1[2] FAD1[3] FAD1[4] FAD1[5] FAD1[6] 
+ FAD1[7] FAD1[8] FAD1[9] FAD1[10] FAD2[0] FAD2[1] FAD2[2] FAD2[3] FAD2[4] 
+ FAD2[5] FAD2[6] FAD2[7] FAD2[8] FAD2[9] FAD2[10] PD PTSEL Q_LL Q_LR REDEN1 
+ REDEN2 RSTB RTSEL[0] RTSEL[1] SCLK SDIN SDOUT TM VDDI VSSI WEB WEBM 
+ WL_TK_ACT[0] WL_TK_ACT[1] WL_TK_ACT[2] WL_TK_ACT[3] WL_TK_ACT[4] 
+ WL_TK_ACT[5] WL_TK_ACT[6] WL_TK_ACT[7] WL_TK_ACT[8] WL_TK_ACT[9] 
+ WL_TK_ACT[10] WL_TK_ACT[11] WL_TK_ACT[12] WL_TK_ACT[13] WL_TK_ACT[14] 
+ WL_TK_ACT[15] WL_TK_ACT[16] WL_TK_ACT[17] WL_TK_ACT[18] WL_TK_ACT[19] 
+ WL_TK_ACT[20] WL_TK_ACT[21] WL_TK_ACT[22] WL_TK_ACT[23] WL_TK_ACT[24] 
+ WL_TK_ACT[25] WL_TK_ACT[26] WL_TK_ACT[27] WL_TK_ACT[28] WL_TK_ACT[29] 
+ WL_TK_ACT[30] WL_TK_ACT[31] WL_TK_ACT[32] WL_TK_ACT[33] WL_TK_ACT[34] 
+ WL_TK_ACT[35] WL_TK_ACT[36] WL_TK_ACT[37] WL_TK_ACT[38] WL_TK_ACT[39] 
+ WL_TK_ACT[40] WL_TK_ACT[41] WL_TK_ACT[42] WL_TK_ACT[43] WL_TK_ACT[44] 
+ WL_TK_ACT[45] WL_TK_ACT[46] WL_TK_ACT[47] WL_TK_ACT[48] WL_TK_ACT[49] 
+ WL_TK_ACT[50] WL_TK_ACT[51] WL_TK_ACT[52] WL_TK_ACT[53] WL_TK_ACT[54] 
+ WL_TK_ACT[55] WL_TK_ACT[56] WL_TK_ACT[57] WL_TK_ACT[58] WL_TK_ACT[59] 
+ WL_TK_ACT[60] WL_TK_ACT[61] WL_TK_ACT[62] WL_TK_ACT[63] WL_TK_ACT[64] 
+ WL_TK_ACT[65] WL_TK_ACT[66] WL_TK_ACT[67] WL_TK_ACT[68] WL_TK_ACT[69] 
+ WL_TK_ACT[70] WL_TK_ACT[71] WL_TK_ACT[72] WL_TK_ACT[73] WL_TK_ACT[74] 
+ WL_TK_ACT[75] WL_TK_ACT[76] WL_TK_ACT[77] WL_TK_ACT[78] WL_TK_ACT[79] 
+ WL_TK_ACT[80] WL_TK_ACT[81] WL_TK_ACT[82] WL_TK_ACT[83] WL_TK_ACT[84] 
+ WL_TK_ACT[85] WL_TK_ACT[86] WL_TK_ACT[87] WL_TK_ACT[88] WL_TK_ACT[89] 
+ WL_TK_ACT[90] WL_TK_ACT[91] WL_TK_ACT[92] WL_TK_ACT[93] WL_TK_ACT[94] 
+ WL_TK_ACT[95] WL_TK_ACT[96] WL_TK_ACT[97] WL_TK_ACT[98] WL_TK_ACT[99] 
+ WL_TK_ACT[100] WL_TK_ACT[101] WL_TK_ACT[102] WL_TK_ACT[103] WL_TK_ACT[104] 
+ WL_TK_ACT[105] WL_TK_ACT[106] WL_TK_ACT[107] WL_TK_ACT[108] WL_TK_ACT[109] 
+ WL_TK_ACT[110] WL_TK_ACT[111] WL_TK_ACT[112] WL_TK_ACT[113] WL_TK_ACT[114] 
+ WL_TK_ACT[115] WL_TK_ACT[116] WL_TK_ACT[117] WL_TK_ACT[118] WL_TK_ACT[119] 
+ WL_TK_ACT[120] WL_TK_ACT[121] WL_TK_ACT[122] WL_TK_ACT[123] WL_TK_ACT[124] 
+ WL_TK_ACT[125] WL_TK_ACT[126] WL_TK_ACT[127] WL_TK_ACT[128] WL_TK_ACT[129] 
+ WL_TK_ACT[130] WL_TK_ACT[131] WL_TK_ACT[132] WL_TK_ACT[133] WL_TK_ACT[134] 
+ WL_TK_ACT[135] WL_TK_ACT[136] WL_TK_ACT[137] WL_TK_ACT[138] WL_TK_ACT[139] 
+ WL_TK_ACT[140] WL_TK_ACT[141] WL_TK_ACT[142] WL_TK_ACT[143] WL_TK_ACT[144] 
+ WL_TK_ACT[145] WL_TK_ACT[146] WL_TK_ACT[147] WL_TK_ACT[148] WL_TK_ACT[149] 
+ WL_TK_ACT[150] WL_TK_ACT[151] WL_TK_ACT[152] WL_TK_ACT[153] WL_TK_ACT[154] 
+ WL_TK_ACT[155] WL_TK_ACT[156] WL_TK_ACT[157] WL_TK_ACT[158] WL_TK_ACT[159] 
+ WL_TK_ACT[160] WL_TK_ACT[161] WL_TK_ACT[162] WL_TK_ACT[163] WL_TK_ACT[164] 
+ WL_TK_ACT[165] WL_TK_ACT[166] WL_TK_ACT[167] WL_TK_ACT[168] WL_TK_ACT[169] 
+ WL_TK_ACT[170] WL_TK_ACT[171] WL_TK_ACT[172] WL_TK_ACT[173] WL_TK_ACT[174] 
+ WL_TK_ACT[175] WL_TK_ACT[176] WL_TK_ACT[177] WL_TK_ACT[178] WL_TK_ACT[179] 
+ WL_TK_ACT[180] WL_TK_ACT[181] WL_TK_ACT[182] WL_TK_ACT[183] WL_TK_ACT[184] 
+ WL_TK_ACT[185] WL_TK_ACT[186] WL_TK_ACT[187] WL_TK_ACT[188] WL_TK_ACT[189] 
+ WL_TK_ACT[190] WL_TK_ACT[191] WL_TK_ACT[192] WL_TK_ACT[193] WL_TK_ACT[194] 
+ WL_TK_ACT[195] WL_TK_ACT[196] WL_TK_ACT[197] WL_TK_ACT[198] WL_TK_ACT[199] 
+ WL_TK_ACT[200] WL_TK_ACT[201] WL_TK_ACT[202] WL_TK_ACT[203] WL_TK_ACT[204] 
+ WL_TK_ACT[205] WL_TK_ACT[206] WL_TK_ACT[207] WL_TK_ACT[208] WL_TK_ACT[209] 
+ WL_TK_ACT[210] WL_TK_ACT[211] WL_TK_ACT[212] WL_TK_ACT[213] WL_TK_ACT[214] 
+ WL_TK_ACT[215] WL_TK_ACT[216] WL_TK_ACT[217] WL_TK_ACT[218] WL_TK_ACT[219] 
+ WL_TK_ACT[220] WL_TK_ACT[221] WL_TK_ACT[222] WL_TK_ACT[223] WL_TK_ACT[224] 
+ WL_TK_ACT[225] WL_TK_ACT[226] WL_TK_ACT[227] WL_TK_ACT[228] WL_TK_ACT[229] 
+ WL_TK_ACT[230] WL_TK_ACT[231] WL_TK_ACT[232] WL_TK_ACT[233] WL_TK_ACT[234] 
+ WL_TK_ACT[235] WL_TK_ACT[236] WL_TK_ACT[237] WL_TK_ACT[238] WL_TK_ACT[239] 
+ WL_TK_ACT[240] WL_TK_ACT[241] WL_TK_ACT[242] WL_TK_ACT[243] WL_TK_ACT[244] 
+ WL_TK_ACT[245] WL_TK_ACT[246] WL_TK_ACT[247] WL_TK_ACT[248] WL_TK_ACT[249] 
+ WL_TK_ACT[250] WL_TK_ACT[251] WL_TK_ACT[252] WL_TK_ACT[253] WL_TK_ACT[254] 
+ WL_TK_ACT[255] WL_TK_ACT[256] WL_TK_ACT[257] WL_TK_ACT[258] WL_TK_ACT[259] 
+ WL_TK_ACT[260] WL_TK_ACT[261] WL_TK_ACT[262] WL_TK_ACT[263] WL_TK_ACT[264] 
+ WL_TK_ACT[265] WL_TK_ACT[266] WL_TK_ACT[267] WL_TK_ACT[268] WL_TK_ACT[269] 
+ WL_TK_ACT[270] WL_TK_ACT[271] WL_TK_ACT[272] WL_TK_ACT[273] WL_TK_ACT[274] 
+ WL_TK_ACT[275] WL_TK_ACT[276] WL_TK_ACT[277] WL_TK_ACT[278] WL_TK_ACT[279] 
+ WL_TK_ACT[280] WL_TK_ACT[281] WL_TK_ACT[282] WL_TK_ACT[283] WL_TK_ACT[284] 
+ WL_TK_ACT[285] WL_TK_ACT[286] WL_TK_ACT[287] WL_TK_ACT[288] WL_TK_ACT[289] 
+ WL_TK_ACT[290] WL_TK_ACT[291] WL_TK_ACT[292] WL_TK_ACT[293] WL_TK_ACT[294] 
+ WL_TK_ACT[295] WL_TK_ACT[296] WL_TK_ACT[297] WL_TK_ACT[298] WL_TK_ACT[299] 
+ WL_TK_ACT[300] WL_TK_ACT[301] WL_TK_ACT[302] WL_TK_ACT[303] WL_TK_ACT[304] 
+ WL_TK_ACT[305] WL_TK_ACT[306] WL_TK_ACT[307] WL_TK_ACT[308] WL_TK_ACT[309] 
+ WL_TK_ACT[310] WL_TK_ACT[311] WL_TK_ACT[312] WL_TK_ACT[313] WL_TK_ACT[314] 
+ WL_TK_ACT[315] WL_TK_ACT[316] WL_TK_ACT[317] WL_TK_ACT[318] WL_TK_ACT[319] 
+ WL_TK_ACT[320] WL_TK_ACT[321] WL_TK_ACT[322] WL_TK_ACT[323] WL_TK_ACT[324] 
+ WL_TK_ACT[325] WL_TK_ACT[326] WL_TK_ACT[327] WL_TK_ACT[328] WL_TK_ACT[329] 
+ WL_TK_ACT[330] WL_TK_ACT[331] WL_TK_ACT[332] WL_TK_ACT[333] WL_TK_ACT[334] 
+ WL_TK_ACT[335] WL_TK_ACT[336] WL_TK_ACT[337] WL_TK_ACT[338] WL_TK_ACT[339] 
+ WL_TK_ACT[340] WL_TK_ACT[341] WL_TK_ACT[342] WL_TK_ACT[343] WL_TK_ACT[344] 
+ WL_TK_ACT[345] WL_TK_ACT[346] WL_TK_ACT[347] WL_TK_ACT[348] WL_TK_ACT[349] 
+ WL_TK_ACT[350] WL_TK_ACT[351] WL_TK_ACT[352] WL_TK_ACT[353] WL_TK_ACT[354] 
+ WL_TK_ACT[355] WL_TK_ACT[356] WL_TK_ACT[357] WL_TK_ACT[358] WL_TK_ACT[359] 
+ WL_TK_ACT[360] WL_TK_ACT[361] WL_TK_ACT[362] WL_TK_ACT[363] WL_TK_ACT[364] 
+ WL_TK_ACT[365] WL_TK_ACT[366] WL_TK_ACT[367] WL_TK_ACT[368] WL_TK_ACT[369] 
+ WL_TK_ACT[370] WL_TK_ACT[371] WL_TK_ACT[372] WL_TK_ACT[373] WL_TK_ACT[374] 
+ WL_TK_ACT[375] WL_TK_ACT[376] WL_TK_ACT[377] WL_TK_ACT[378] WL_TK_ACT[379] 
+ WL_TK_ACT[380] WL_TK_ACT[381] WL_TK_ACT[382] WL_TK_ACT[383] WL_TK_ACT[384] 
+ WL_TK_ACT[385] WL_TK_ACT[386] WL_TK_ACT[387] WL_TK_ACT[388] WL_TK_ACT[389] 
+ WL_TK_ACT[390] WL_TK_ACT[391] WL_TK_ACT[392] WL_TK_ACT[393] WL_TK_ACT[394] 
+ WL_TK_ACT[395] WL_TK_ACT[396] WL_TK_ACT[397] WL_TK_ACT[398] WL_TK_ACT[399] 
+ WL_TK_ACT[400] WL_TK_ACT[401] WL_TK_ACT[402] WL_TK_ACT[403] WL_TK_ACT[404] 
+ WL_TK_ACT[405] WL_TK_ACT[406] WL_TK_ACT[407] WL_TK_ACT[408] WL_TK_ACT[409] 
+ WL_TK_ACT[410] WL_TK_ACT[411] WL_TK_ACT[412] WL_TK_ACT[413] WL_TK_ACT[414] 
+ WL_TK_ACT[415] WL_TK_ACT[416] WL_TK_ACT[417] WL_TK_ACT[418] WL_TK_ACT[419] 
+ WL_TK_ACT[420] WL_TK_ACT[421] WL_TK_ACT[422] WL_TK_ACT[423] WL_TK_ACT[424] 
+ WL_TK_ACT[425] WL_TK_ACT[426] WL_TK_ACT[427] WL_TK_ACT[428] WL_TK_ACT[429] 
+ WL_TK_ACT[430] WL_TK_ACT[431] WL_TK_ACT[432] WL_TK_ACT[433] WL_TK_ACT[434] 
+ WL_TK_ACT[435] WL_TK_ACT[436] WL_TK_ACT[437] WL_TK_ACT[438] WL_TK_ACT[439] 
+ WL_TK_ACT[440] WL_TK_ACT[441] WL_TK_ACT[442] WL_TK_ACT[443] WL_TK_ACT[444] 
+ WL_TK_ACT[445] WL_TK_ACT[446] WL_TK_ACT[447] WL_TK_ACT[448] WL_TK_ACT[449] 
+ WL_TK_ACT[450] WL_TK_ACT[451] WL_TK_ACT[452] WL_TK_ACT[453] WL_TK_ACT[454] 
+ WL_TK_ACT[455] WL_TK_ACT[456] WL_TK_ACT[457] WL_TK_ACT[458] WL_TK_ACT[459] 
+ WL_TK_ACT[460] WL_TK_ACT[461] WL_TK_ACT[462] WL_TK_ACT[463] WL_TK_ACT[464] 
+ WL_TK_ACT[465] WL_TK_ACT[466] WL_TK_ACT[467] WL_TK_ACT[468] WL_TK_ACT[469] 
+ WL_TK_ACT[470] WL_TK_ACT[471] WL_TK_ACT[472] WL_TK_ACT[473] WL_TK_ACT[474] 
+ WL_TK_ACT[475] WL_TK_ACT[476] WL_TK_ACT[477] WL_TK_ACT[478] WL_TK_ACT[479] 
+ WL_TK_ACT[480] WL_TK_ACT[481] WL_TK_ACT[482] WL_TK_ACT[483] WL_TK_ACT[484] 
+ WL_TK_ACT[485] WL_TK_ACT[486] WL_TK_ACT[487] WL_TK_ACT[488] WL_TK_ACT[489] 
+ WL_TK_ACT[490] WL_TK_ACT[491] WL_TK_ACT[492] WL_TK_ACT[493] WL_TK_ACT[494] 
+ WL_TK_ACT[495] WL_TK_ACT[496] WL_TK_ACT[497] WL_TK_ACT[498] WL_TK_ACT[499] 
+ WL_TK_ACT[500] WL_TK_ACT[501] WL_TK_ACT[502] WL_TK_ACT[503] WL_TK_ACT[504] 
+ WL_TK_ACT[505] WL_TK_ACT[506] WL_TK_ACT[507] WL_TK_ACT[508] WL_TK_ACT[509] 
+ WL_TK_ACT[510] WL_TK_ACT[511] WL_TK_LD WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] 
+ X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] 
+ XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YM[0] YM[1] YM[2] 
+ YM[3]
*.PININFO AWT:I BIST:I BWEBM_LL:I BWEBM_LR:I BWEB_LL:I BWEB_LR:I CEB:I CEBM:I 
*.PININFO CLK:I DM_LL:I DM_LR:I D_LL:I D_LR:I FAD1[0]:I FAD1[1]:I FAD1[2]:I 
*.PININFO FAD1[3]:I FAD1[4]:I FAD1[5]:I FAD1[6]:I FAD1[7]:I FAD1[8]:I 
*.PININFO FAD1[9]:I FAD1[10]:I FAD2[0]:I FAD2[1]:I FAD2[2]:I FAD2[3]:I 
*.PININFO FAD2[4]:I FAD2[5]:I FAD2[6]:I FAD2[7]:I FAD2[8]:I FAD2[9]:I 
*.PININFO FAD2[10]:I PD:I PTSEL:I REDEN1:I REDEN2:I RSTB:I RTSEL[0]:I 
*.PININFO RTSEL[1]:I SCLK:I SDIN:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I 
*.PININFO XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I 
*.PININFO Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I Q_LL:O Q_LR:O SDOUT:O 
*.PININFO VDDI:B VSSI:B WL_TK_ACT[0]:B WL_TK_ACT[1]:B WL_TK_ACT[2]:B 
*.PININFO WL_TK_ACT[3]:B WL_TK_ACT[4]:B WL_TK_ACT[5]:B WL_TK_ACT[6]:B 
*.PININFO WL_TK_ACT[7]:B WL_TK_ACT[8]:B WL_TK_ACT[9]:B WL_TK_ACT[10]:B 
*.PININFO WL_TK_ACT[11]:B WL_TK_ACT[12]:B WL_TK_ACT[13]:B WL_TK_ACT[14]:B 
*.PININFO WL_TK_ACT[15]:B WL_TK_ACT[16]:B WL_TK_ACT[17]:B WL_TK_ACT[18]:B 
*.PININFO WL_TK_ACT[19]:B WL_TK_ACT[20]:B WL_TK_ACT[21]:B WL_TK_ACT[22]:B 
*.PININFO WL_TK_ACT[23]:B WL_TK_ACT[24]:B WL_TK_ACT[25]:B WL_TK_ACT[26]:B 
*.PININFO WL_TK_ACT[27]:B WL_TK_ACT[28]:B WL_TK_ACT[29]:B WL_TK_ACT[30]:B 
*.PININFO WL_TK_ACT[31]:B WL_TK_ACT[32]:B WL_TK_ACT[33]:B WL_TK_ACT[34]:B 
*.PININFO WL_TK_ACT[35]:B WL_TK_ACT[36]:B WL_TK_ACT[37]:B WL_TK_ACT[38]:B 
*.PININFO WL_TK_ACT[39]:B WL_TK_ACT[40]:B WL_TK_ACT[41]:B WL_TK_ACT[42]:B 
*.PININFO WL_TK_ACT[43]:B WL_TK_ACT[44]:B WL_TK_ACT[45]:B WL_TK_ACT[46]:B 
*.PININFO WL_TK_ACT[47]:B WL_TK_ACT[48]:B WL_TK_ACT[49]:B WL_TK_ACT[50]:B 
*.PININFO WL_TK_ACT[51]:B WL_TK_ACT[52]:B WL_TK_ACT[53]:B WL_TK_ACT[54]:B 
*.PININFO WL_TK_ACT[55]:B WL_TK_ACT[56]:B WL_TK_ACT[57]:B WL_TK_ACT[58]:B 
*.PININFO WL_TK_ACT[59]:B WL_TK_ACT[60]:B WL_TK_ACT[61]:B WL_TK_ACT[62]:B 
*.PININFO WL_TK_ACT[63]:B WL_TK_ACT[64]:B WL_TK_ACT[65]:B WL_TK_ACT[66]:B 
*.PININFO WL_TK_ACT[67]:B WL_TK_ACT[68]:B WL_TK_ACT[69]:B WL_TK_ACT[70]:B 
*.PININFO WL_TK_ACT[71]:B WL_TK_ACT[72]:B WL_TK_ACT[73]:B WL_TK_ACT[74]:B 
*.PININFO WL_TK_ACT[75]:B WL_TK_ACT[76]:B WL_TK_ACT[77]:B WL_TK_ACT[78]:B 
*.PININFO WL_TK_ACT[79]:B WL_TK_ACT[80]:B WL_TK_ACT[81]:B WL_TK_ACT[82]:B 
*.PININFO WL_TK_ACT[83]:B WL_TK_ACT[84]:B WL_TK_ACT[85]:B WL_TK_ACT[86]:B 
*.PININFO WL_TK_ACT[87]:B WL_TK_ACT[88]:B WL_TK_ACT[89]:B WL_TK_ACT[90]:B 
*.PININFO WL_TK_ACT[91]:B WL_TK_ACT[92]:B WL_TK_ACT[93]:B WL_TK_ACT[94]:B 
*.PININFO WL_TK_ACT[95]:B WL_TK_ACT[96]:B WL_TK_ACT[97]:B WL_TK_ACT[98]:B 
*.PININFO WL_TK_ACT[99]:B WL_TK_ACT[100]:B WL_TK_ACT[101]:B WL_TK_ACT[102]:B 
*.PININFO WL_TK_ACT[103]:B WL_TK_ACT[104]:B WL_TK_ACT[105]:B WL_TK_ACT[106]:B 
*.PININFO WL_TK_ACT[107]:B WL_TK_ACT[108]:B WL_TK_ACT[109]:B WL_TK_ACT[110]:B 
*.PININFO WL_TK_ACT[111]:B WL_TK_ACT[112]:B WL_TK_ACT[113]:B WL_TK_ACT[114]:B 
*.PININFO WL_TK_ACT[115]:B WL_TK_ACT[116]:B WL_TK_ACT[117]:B WL_TK_ACT[118]:B 
*.PININFO WL_TK_ACT[119]:B WL_TK_ACT[120]:B WL_TK_ACT[121]:B WL_TK_ACT[122]:B 
*.PININFO WL_TK_ACT[123]:B WL_TK_ACT[124]:B WL_TK_ACT[125]:B WL_TK_ACT[126]:B 
*.PININFO WL_TK_ACT[127]:B WL_TK_ACT[128]:B WL_TK_ACT[129]:B WL_TK_ACT[130]:B 
*.PININFO WL_TK_ACT[131]:B WL_TK_ACT[132]:B WL_TK_ACT[133]:B WL_TK_ACT[134]:B 
*.PININFO WL_TK_ACT[135]:B WL_TK_ACT[136]:B WL_TK_ACT[137]:B WL_TK_ACT[138]:B 
*.PININFO WL_TK_ACT[139]:B WL_TK_ACT[140]:B WL_TK_ACT[141]:B WL_TK_ACT[142]:B 
*.PININFO WL_TK_ACT[143]:B WL_TK_ACT[144]:B WL_TK_ACT[145]:B WL_TK_ACT[146]:B 
*.PININFO WL_TK_ACT[147]:B WL_TK_ACT[148]:B WL_TK_ACT[149]:B WL_TK_ACT[150]:B 
*.PININFO WL_TK_ACT[151]:B WL_TK_ACT[152]:B WL_TK_ACT[153]:B WL_TK_ACT[154]:B 
*.PININFO WL_TK_ACT[155]:B WL_TK_ACT[156]:B WL_TK_ACT[157]:B WL_TK_ACT[158]:B 
*.PININFO WL_TK_ACT[159]:B WL_TK_ACT[160]:B WL_TK_ACT[161]:B WL_TK_ACT[162]:B 
*.PININFO WL_TK_ACT[163]:B WL_TK_ACT[164]:B WL_TK_ACT[165]:B WL_TK_ACT[166]:B 
*.PININFO WL_TK_ACT[167]:B WL_TK_ACT[168]:B WL_TK_ACT[169]:B WL_TK_ACT[170]:B 
*.PININFO WL_TK_ACT[171]:B WL_TK_ACT[172]:B WL_TK_ACT[173]:B WL_TK_ACT[174]:B 
*.PININFO WL_TK_ACT[175]:B WL_TK_ACT[176]:B WL_TK_ACT[177]:B WL_TK_ACT[178]:B 
*.PININFO WL_TK_ACT[179]:B WL_TK_ACT[180]:B WL_TK_ACT[181]:B WL_TK_ACT[182]:B 
*.PININFO WL_TK_ACT[183]:B WL_TK_ACT[184]:B WL_TK_ACT[185]:B WL_TK_ACT[186]:B 
*.PININFO WL_TK_ACT[187]:B WL_TK_ACT[188]:B WL_TK_ACT[189]:B WL_TK_ACT[190]:B 
*.PININFO WL_TK_ACT[191]:B WL_TK_ACT[192]:B WL_TK_ACT[193]:B WL_TK_ACT[194]:B 
*.PININFO WL_TK_ACT[195]:B WL_TK_ACT[196]:B WL_TK_ACT[197]:B WL_TK_ACT[198]:B 
*.PININFO WL_TK_ACT[199]:B WL_TK_ACT[200]:B WL_TK_ACT[201]:B WL_TK_ACT[202]:B 
*.PININFO WL_TK_ACT[203]:B WL_TK_ACT[204]:B WL_TK_ACT[205]:B WL_TK_ACT[206]:B 
*.PININFO WL_TK_ACT[207]:B WL_TK_ACT[208]:B WL_TK_ACT[209]:B WL_TK_ACT[210]:B 
*.PININFO WL_TK_ACT[211]:B WL_TK_ACT[212]:B WL_TK_ACT[213]:B WL_TK_ACT[214]:B 
*.PININFO WL_TK_ACT[215]:B WL_TK_ACT[216]:B WL_TK_ACT[217]:B WL_TK_ACT[218]:B 
*.PININFO WL_TK_ACT[219]:B WL_TK_ACT[220]:B WL_TK_ACT[221]:B WL_TK_ACT[222]:B 
*.PININFO WL_TK_ACT[223]:B WL_TK_ACT[224]:B WL_TK_ACT[225]:B WL_TK_ACT[226]:B 
*.PININFO WL_TK_ACT[227]:B WL_TK_ACT[228]:B WL_TK_ACT[229]:B WL_TK_ACT[230]:B 
*.PININFO WL_TK_ACT[231]:B WL_TK_ACT[232]:B WL_TK_ACT[233]:B WL_TK_ACT[234]:B 
*.PININFO WL_TK_ACT[235]:B WL_TK_ACT[236]:B WL_TK_ACT[237]:B WL_TK_ACT[238]:B 
*.PININFO WL_TK_ACT[239]:B WL_TK_ACT[240]:B WL_TK_ACT[241]:B WL_TK_ACT[242]:B 
*.PININFO WL_TK_ACT[243]:B WL_TK_ACT[244]:B WL_TK_ACT[245]:B WL_TK_ACT[246]:B 
*.PININFO WL_TK_ACT[247]:B WL_TK_ACT[248]:B WL_TK_ACT[249]:B WL_TK_ACT[250]:B 
*.PININFO WL_TK_ACT[251]:B WL_TK_ACT[252]:B WL_TK_ACT[253]:B WL_TK_ACT[254]:B 
*.PININFO WL_TK_ACT[255]:B WL_TK_ACT[256]:B WL_TK_ACT[257]:B WL_TK_ACT[258]:B 
*.PININFO WL_TK_ACT[259]:B WL_TK_ACT[260]:B WL_TK_ACT[261]:B WL_TK_ACT[262]:B 
*.PININFO WL_TK_ACT[263]:B WL_TK_ACT[264]:B WL_TK_ACT[265]:B WL_TK_ACT[266]:B 
*.PININFO WL_TK_ACT[267]:B WL_TK_ACT[268]:B WL_TK_ACT[269]:B WL_TK_ACT[270]:B 
*.PININFO WL_TK_ACT[271]:B WL_TK_ACT[272]:B WL_TK_ACT[273]:B WL_TK_ACT[274]:B 
*.PININFO WL_TK_ACT[275]:B WL_TK_ACT[276]:B WL_TK_ACT[277]:B WL_TK_ACT[278]:B 
*.PININFO WL_TK_ACT[279]:B WL_TK_ACT[280]:B WL_TK_ACT[281]:B WL_TK_ACT[282]:B 
*.PININFO WL_TK_ACT[283]:B WL_TK_ACT[284]:B WL_TK_ACT[285]:B WL_TK_ACT[286]:B 
*.PININFO WL_TK_ACT[287]:B WL_TK_ACT[288]:B WL_TK_ACT[289]:B WL_TK_ACT[290]:B 
*.PININFO WL_TK_ACT[291]:B WL_TK_ACT[292]:B WL_TK_ACT[293]:B WL_TK_ACT[294]:B 
*.PININFO WL_TK_ACT[295]:B WL_TK_ACT[296]:B WL_TK_ACT[297]:B WL_TK_ACT[298]:B 
*.PININFO WL_TK_ACT[299]:B WL_TK_ACT[300]:B WL_TK_ACT[301]:B WL_TK_ACT[302]:B 
*.PININFO WL_TK_ACT[303]:B WL_TK_ACT[304]:B WL_TK_ACT[305]:B WL_TK_ACT[306]:B 
*.PININFO WL_TK_ACT[307]:B WL_TK_ACT[308]:B WL_TK_ACT[309]:B WL_TK_ACT[310]:B 
*.PININFO WL_TK_ACT[311]:B WL_TK_ACT[312]:B WL_TK_ACT[313]:B WL_TK_ACT[314]:B 
*.PININFO WL_TK_ACT[315]:B WL_TK_ACT[316]:B WL_TK_ACT[317]:B WL_TK_ACT[318]:B 
*.PININFO WL_TK_ACT[319]:B WL_TK_ACT[320]:B WL_TK_ACT[321]:B WL_TK_ACT[322]:B 
*.PININFO WL_TK_ACT[323]:B WL_TK_ACT[324]:B WL_TK_ACT[325]:B WL_TK_ACT[326]:B 
*.PININFO WL_TK_ACT[327]:B WL_TK_ACT[328]:B WL_TK_ACT[329]:B WL_TK_ACT[330]:B 
*.PININFO WL_TK_ACT[331]:B WL_TK_ACT[332]:B WL_TK_ACT[333]:B WL_TK_ACT[334]:B 
*.PININFO WL_TK_ACT[335]:B WL_TK_ACT[336]:B WL_TK_ACT[337]:B WL_TK_ACT[338]:B 
*.PININFO WL_TK_ACT[339]:B WL_TK_ACT[340]:B WL_TK_ACT[341]:B WL_TK_ACT[342]:B 
*.PININFO WL_TK_ACT[343]:B WL_TK_ACT[344]:B WL_TK_ACT[345]:B WL_TK_ACT[346]:B 
*.PININFO WL_TK_ACT[347]:B WL_TK_ACT[348]:B WL_TK_ACT[349]:B WL_TK_ACT[350]:B 
*.PININFO WL_TK_ACT[351]:B WL_TK_ACT[352]:B WL_TK_ACT[353]:B WL_TK_ACT[354]:B 
*.PININFO WL_TK_ACT[355]:B WL_TK_ACT[356]:B WL_TK_ACT[357]:B WL_TK_ACT[358]:B 
*.PININFO WL_TK_ACT[359]:B WL_TK_ACT[360]:B WL_TK_ACT[361]:B WL_TK_ACT[362]:B 
*.PININFO WL_TK_ACT[363]:B WL_TK_ACT[364]:B WL_TK_ACT[365]:B WL_TK_ACT[366]:B 
*.PININFO WL_TK_ACT[367]:B WL_TK_ACT[368]:B WL_TK_ACT[369]:B WL_TK_ACT[370]:B 
*.PININFO WL_TK_ACT[371]:B WL_TK_ACT[372]:B WL_TK_ACT[373]:B WL_TK_ACT[374]:B 
*.PININFO WL_TK_ACT[375]:B WL_TK_ACT[376]:B WL_TK_ACT[377]:B WL_TK_ACT[378]:B 
*.PININFO WL_TK_ACT[379]:B WL_TK_ACT[380]:B WL_TK_ACT[381]:B WL_TK_ACT[382]:B 
*.PININFO WL_TK_ACT[383]:B WL_TK_ACT[384]:B WL_TK_ACT[385]:B WL_TK_ACT[386]:B 
*.PININFO WL_TK_ACT[387]:B WL_TK_ACT[388]:B WL_TK_ACT[389]:B WL_TK_ACT[390]:B 
*.PININFO WL_TK_ACT[391]:B WL_TK_ACT[392]:B WL_TK_ACT[393]:B WL_TK_ACT[394]:B 
*.PININFO WL_TK_ACT[395]:B WL_TK_ACT[396]:B WL_TK_ACT[397]:B WL_TK_ACT[398]:B 
*.PININFO WL_TK_ACT[399]:B WL_TK_ACT[400]:B WL_TK_ACT[401]:B WL_TK_ACT[402]:B 
*.PININFO WL_TK_ACT[403]:B WL_TK_ACT[404]:B WL_TK_ACT[405]:B WL_TK_ACT[406]:B 
*.PININFO WL_TK_ACT[407]:B WL_TK_ACT[408]:B WL_TK_ACT[409]:B WL_TK_ACT[410]:B 
*.PININFO WL_TK_ACT[411]:B WL_TK_ACT[412]:B WL_TK_ACT[413]:B WL_TK_ACT[414]:B 
*.PININFO WL_TK_ACT[415]:B WL_TK_ACT[416]:B WL_TK_ACT[417]:B WL_TK_ACT[418]:B 
*.PININFO WL_TK_ACT[419]:B WL_TK_ACT[420]:B WL_TK_ACT[421]:B WL_TK_ACT[422]:B 
*.PININFO WL_TK_ACT[423]:B WL_TK_ACT[424]:B WL_TK_ACT[425]:B WL_TK_ACT[426]:B 
*.PININFO WL_TK_ACT[427]:B WL_TK_ACT[428]:B WL_TK_ACT[429]:B WL_TK_ACT[430]:B 
*.PININFO WL_TK_ACT[431]:B WL_TK_ACT[432]:B WL_TK_ACT[433]:B WL_TK_ACT[434]:B 
*.PININFO WL_TK_ACT[435]:B WL_TK_ACT[436]:B WL_TK_ACT[437]:B WL_TK_ACT[438]:B 
*.PININFO WL_TK_ACT[439]:B WL_TK_ACT[440]:B WL_TK_ACT[441]:B WL_TK_ACT[442]:B 
*.PININFO WL_TK_ACT[443]:B WL_TK_ACT[444]:B WL_TK_ACT[445]:B WL_TK_ACT[446]:B 
*.PININFO WL_TK_ACT[447]:B WL_TK_ACT[448]:B WL_TK_ACT[449]:B WL_TK_ACT[450]:B 
*.PININFO WL_TK_ACT[451]:B WL_TK_ACT[452]:B WL_TK_ACT[453]:B WL_TK_ACT[454]:B 
*.PININFO WL_TK_ACT[455]:B WL_TK_ACT[456]:B WL_TK_ACT[457]:B WL_TK_ACT[458]:B 
*.PININFO WL_TK_ACT[459]:B WL_TK_ACT[460]:B WL_TK_ACT[461]:B WL_TK_ACT[462]:B 
*.PININFO WL_TK_ACT[463]:B WL_TK_ACT[464]:B WL_TK_ACT[465]:B WL_TK_ACT[466]:B 
*.PININFO WL_TK_ACT[467]:B WL_TK_ACT[468]:B WL_TK_ACT[469]:B WL_TK_ACT[470]:B 
*.PININFO WL_TK_ACT[471]:B WL_TK_ACT[472]:B WL_TK_ACT[473]:B WL_TK_ACT[474]:B 
*.PININFO WL_TK_ACT[475]:B WL_TK_ACT[476]:B WL_TK_ACT[477]:B WL_TK_ACT[478]:B 
*.PININFO WL_TK_ACT[479]:B WL_TK_ACT[480]:B WL_TK_ACT[481]:B WL_TK_ACT[482]:B 
*.PININFO WL_TK_ACT[483]:B WL_TK_ACT[484]:B WL_TK_ACT[485]:B WL_TK_ACT[486]:B 
*.PININFO WL_TK_ACT[487]:B WL_TK_ACT[488]:B WL_TK_ACT[489]:B WL_TK_ACT[490]:B 
*.PININFO WL_TK_ACT[491]:B WL_TK_ACT[492]:B WL_TK_ACT[493]:B WL_TK_ACT[494]:B 
*.PININFO WL_TK_ACT[495]:B WL_TK_ACT[496]:B WL_TK_ACT[497]:B WL_TK_ACT[498]:B 
*.PININFO WL_TK_ACT[499]:B WL_TK_ACT[500]:B WL_TK_ACT[501]:B WL_TK_ACT[502]:B 
*.PININFO WL_TK_ACT[503]:B WL_TK_ACT[504]:B WL_TK_ACT[505]:B WL_TK_ACT[506]:B 
*.PININFO WL_TK_ACT[507]:B WL_TK_ACT[508]:B WL_TK_ACT[509]:B WL_TK_ACT[510]:B 
*.PININFO WL_TK_ACT[511]:B WL_TK_LD:B
XBK_WLDV_U VDDHD VDDI DEC_X0_7[0] DEC_X0_7[1] DEC_X0_7[2] DEC_X0_7[3] 
+ DEC_X0_7[4] DEC_X0_7[5] DEC_X0_7[6] DEC_X0_7[7] NET01202[0] NET01202[1] 
+ NET01202[2] NET01202[3] NET01202[4] NET01202[5] NET01202[6] NET01202[7] 
+ DEC_X1_7[0] DEC_X1_7[1] DEC_X1_7[2] DEC_X1_7[3] DEC_X1_7[4] DEC_X1_7[5] 
+ DEC_X1_7[6] DEC_X1_7[7] NET050[0] NET050[1] NET050[2] NET050[3] NET050[4] 
+ NET050[5] NET050[6] NET050[7] DEC_X2_7[0] DEC_X2_7[1] DEC_X2_7[2] 
+ DEC_X2_7[3] NET051[0] NET051[1] NET051[2] NET051[3] DEC_X3_7[0] DEC_X3_7[1] 
+ DEC_X3_7[2] DEC_X3_7[3] DEC_X3_7[4] DEC_X3_7[5] DEC_X3_7[6] DEC_X3_7[7] 
+ NET01205[0] NET01205[1] NET01205[2] NET01205[3] NET01205[4] NET01205[5] 
+ NET01205[6] NET01205[7] DEC_Y_7[0] DEC_Y_7[1] DEC_Y_7[2] DEC_Y_7[3] 
+ DEC_Y_7[4] DEC_Y_7[5] DEC_Y_7[6] DEC_Y_7[7] NET01201[0] NET01201[1] 
+ NET01201[2] NET01201[3] NET01201[4] NET01201[5] NET01201[6] NET01201[7] 
+ PD_BUF_7 NET01203 PD_CVDDBUF_7 NET01204 RW_RE_7 NET052 VDDHD VDDI VSSI 
+ WLPYB_7 NET1176 WLPY_7 NET1209 WLP_SAE_7 WLP_SAE_TK_7 WLP_SAE_TK_8 WLP_SAE_8 
+ WL_LU1[0] WL_LU1[1] WL_RU1[0] WL_RU1[1] YL_7[0] NET01200 S1AHSF400W40_BK_WLDV_U_SIM
XBK_WLDV_D VDDHD VDDI DEC_X0_1[0] DEC_X0_1[1] DEC_X0_1[2] DEC_X0_1[3] 
+ DEC_X0_1[4] DEC_X0_1[5] DEC_X0_1[6] DEC_X0_1[7] DEC_X0_2[0] DEC_X0_2[1] 
+ DEC_X0_2[2] DEC_X0_2[3] DEC_X0_2[4] DEC_X0_2[5] DEC_X0_2[6] DEC_X0_2[7] 
+ DEC_X1_1[0] DEC_X1_1[1] DEC_X1_1[2] DEC_X1_1[3] DEC_X1_1[4] DEC_X1_1[5] 
+ DEC_X1_1[6] DEC_X1_1[7] DEC_X1_2[0] DEC_X1_2[1] DEC_X1_2[2] DEC_X1_2[3] 
+ DEC_X1_2[4] DEC_X1_2[5] DEC_X1_2[6] DEC_X1_2[7] DEC_X2_1[0] DEC_X2_1[1] 
+ DEC_X2_1[2] DEC_X2_1[3] DEC_X2_2[0] DEC_X2_2[1] DEC_X2_2[2] DEC_X2_2[3] 
+ DEC_X3_1[0] DEC_X3_1[1] DEC_X3_1[2] DEC_X3_1[3] DEC_X3_1[4] DEC_X3_1[5] 
+ DEC_X3_1[6] DEC_X3_1[7] DEC_X3_2[0] DEC_X3_2[1] DEC_X3_2[2] DEC_X3_2[3] 
+ DEC_X3_2[4] DEC_X3_2[5] DEC_X3_2[6] DEC_X3_2[7] DEC_Y_1[0] DEC_Y_1[1] 
+ DEC_Y_1[2] DEC_Y_1[3] DEC_Y_1[4] DEC_Y_1[5] DEC_Y_1[6] DEC_Y_1[7] DEC_Y_2[0] 
+ DEC_Y_2[1] DEC_Y_2[2] DEC_Y_2[3] DEC_Y_2[4] DEC_Y_2[5] DEC_Y_2[6] DEC_Y_2[7] 
+ PD_BUF_1 PD_BUF_2 PD_CVDDBUF_1 PD_CVDDBUF_2 RW_RE_1 RW_RE_2 VDDHD VDDI VSSI 
+ NET129 WLPYB_2 NET130 WLPY_2 WLP_SAE_1 WLP_SAE_TK_1 WLP_SAE_TK_2 WLP_SAE_2 
+ WL_LD1[0] WL_LD1[1] WL_RD1[0] WL_RD1[1] YL_1[0] YL_2[0] S1AHSF400W40_BK_WLDV_D_SIM
XWLPY_LD_U VDDHD VDDI VDDHD VDDI VSSI WLPYB_6 WLPYB_7 WLPY_6 WLPY_7 
+ S1AHSF400W40_WLPY_LD_SIM
XWLPY_LD_D VDDHD VDDI VDDHD VDDI VSSI WLPYB_2 WLPYB_3 WLPY_2 WLPY_3 
+ S1AHSF400W40_WLPY_LD_SIM
XBK_LCNT_D BLEQ_DN_LD1 BLEQ_DN_RD1 BLEQ_UP_LD1 BLEQ_UP_RD1 VDDHD VDDI 
+ DEC_X0_3[0] DEC_X0_3[1] DEC_X0_3[2] DEC_X0_3[3] DEC_X0_3[4] DEC_X0_3[5] 
+ DEC_X0_3[6] DEC_X0_3[7] DEC_X0_4[0] DEC_X0_4[1] DEC_X0_4[2] DEC_X0_4[3] 
+ DEC_X0_4[4] DEC_X0_4[5] DEC_X0_4[6] DEC_X0_4[7] DEC_X1_3[0] DEC_X1_3[1] 
+ DEC_X1_3[2] DEC_X1_3[3] DEC_X1_3[4] DEC_X1_3[5] DEC_X1_3[6] DEC_X1_3[7] 
+ DEC_X1_4[0] DEC_X1_4[1] DEC_X1_4[2] DEC_X1_4[3] DEC_X1_4[4] DEC_X1_4[5] 
+ DEC_X1_4[6] DEC_X1_4[7] DEC_X2_3[0] DEC_X2_3[1] DEC_X2_3[2] DEC_X2_3[3] 
+ DEC_X2_4[0] DEC_X2_4[1] DEC_X2_4[2] DEC_X2_4[3] DEC_X3_3[0] DEC_X3_3[1] 
+ DEC_X3_3[2] DEC_X3_3[3] DEC_X3_3[4] DEC_X3_3[5] DEC_X3_3[6] DEC_X3_3[7] 
+ DEC_X3_4[0] DEC_X3_4[1] DEC_X3_4[2] DEC_X3_4[3] DEC_X3_4[4] DEC_X3_4[5] 
+ DEC_X3_4[6] DEC_X3_4[7] DEC_Y_3[0] DEC_Y_3[1] DEC_Y_3[2] DEC_Y_3[3] 
+ DEC_Y_3[4] DEC_Y_3[5] DEC_Y_3[6] DEC_Y_3[7] Y_DN_LD1[0] Y_DN_LD1[1] 
+ Y_DN_LD1[2] Y_DN_LD1[3] Y_DN_LD1[4] Y_DN_LD1[5] Y_DN_LD1[6] Y_DN_LD1[7] 
+ Y_DN_RD1[0] Y_DN_RD1[1] Y_DN_RD1[2] Y_DN_RD1[3] Y_DN_RD1[4] Y_DN_RD1[5] 
+ Y_DN_RD1[6] Y_DN_RD1[7] DEC_Y_4[0] DEC_Y_4[1] DEC_Y_4[2] DEC_Y_4[3] 
+ DEC_Y_4[4] DEC_Y_4[5] DEC_Y_4[6] DEC_Y_4[7] Y_UP_LD1[0] Y_UP_LD1[1] 
+ Y_UP_LD1[2] Y_UP_LD1[3] Y_UP_LD1[4] Y_UP_LD1[5] Y_UP_LD1[6] Y_UP_LD1[7] 
+ Y_UP_RD1[0] Y_UP_RD1[1] Y_UP_RD1[2] Y_UP_RD1[3] Y_UP_RD1[4] Y_UP_RD1[5] 
+ Y_UP_RD1[6] Y_UP_RD1[7] PD_BUF_3 PD_BUF_4 PD_CVDDBUF_3 PD_CVDDBUF_4 RE_LD1 
+ RE_RD1 RW_RE_3 RW_RE_4 SAEB_LD1 SAEB_RD1 VDDHD VDDI VSSI WE_LD1 WE_RD1 
+ WLPYB_3 NET180 WLPY_3 NET178 WLP_SAE_3 WLP_SAE_TK_3 WLP_SAE_TK_4 WLP_SAE_4 
+ YL_3[0] YL_LD1[0] YL_LD1[1] YL_RD1[0] YL_RD1[1] YL_4[0] S1AHSF400W40_BK_LCNT_D_SIM
XBK_LCNT_U BLEQ_DN_LU1 BLEQ_DN_RU1 BLEQ_UP_LU1 BLEQ_UP_RU1 VDDHD VDDI 
+ DEC_X0_5[0] DEC_X0_5[1] DEC_X0_5[2] DEC_X0_5[3] DEC_X0_5[4] DEC_X0_5[5] 
+ DEC_X0_5[6] DEC_X0_5[7] DEC_X0_6[0] DEC_X0_6[1] DEC_X0_6[2] DEC_X0_6[3] 
+ DEC_X0_6[4] DEC_X0_6[5] DEC_X0_6[6] DEC_X0_6[7] DEC_X1_5[0] DEC_X1_5[1] 
+ DEC_X1_5[2] DEC_X1_5[3] DEC_X1_5[4] DEC_X1_5[5] DEC_X1_5[6] DEC_X1_5[7] 
+ DEC_X1_6[0] DEC_X1_6[1] DEC_X1_6[2] DEC_X1_6[3] DEC_X1_6[4] DEC_X1_6[5] 
+ DEC_X1_6[6] DEC_X1_6[7] DEC_X2_5[0] DEC_X2_5[1] DEC_X2_5[2] DEC_X2_5[3] 
+ DEC_X2_6[0] DEC_X2_6[1] DEC_X2_6[2] DEC_X2_6[3] DEC_X3_5[0] DEC_X3_5[1] 
+ DEC_X3_5[2] DEC_X3_5[3] DEC_X3_5[4] DEC_X3_5[5] DEC_X3_5[6] DEC_X3_5[7] 
+ DEC_X3_6[0] DEC_X3_6[1] DEC_X3_6[2] DEC_X3_6[3] DEC_X3_6[4] DEC_X3_6[5] 
+ DEC_X3_6[6] DEC_X3_6[7] DEC_Y_5[0] DEC_Y_5[1] DEC_Y_5[2] DEC_Y_5[3] 
+ DEC_Y_5[4] DEC_Y_5[5] DEC_Y_5[6] DEC_Y_5[7] Y_DN_LU1[0] Y_DN_LU1[1] 
+ Y_DN_LU1[2] Y_DN_LU1[3] Y_DN_LU1[4] Y_DN_LU1[5] Y_DN_LU1[6] Y_DN_LU1[7] 
+ Y_DN_RU1[0] Y_DN_RU1[1] Y_DN_RU1[2] Y_DN_RU1[3] Y_DN_RU1[4] Y_DN_RU1[5] 
+ Y_DN_RU1[6] Y_DN_RU1[7] DEC_Y_6[0] DEC_Y_6[1] DEC_Y_6[2] DEC_Y_6[3] 
+ DEC_Y_6[4] DEC_Y_6[5] DEC_Y_6[6] DEC_Y_6[7] Y_UP_LU1[0] Y_UP_LU1[1] 
+ Y_UP_LU1[2] Y_UP_LU1[3] Y_UP_LU1[4] Y_UP_LU1[5] Y_UP_LU1[6] Y_UP_LU1[7] 
+ Y_UP_RU1[0] Y_UP_RU1[1] Y_UP_RU1[2] Y_UP_RU1[3] Y_UP_RU1[4] Y_UP_RU1[5] 
+ Y_UP_RU1[6] Y_UP_RU1[7] PD_BUF_5 PD_BUF_6 PD_CVDDBUF_5 PD_CVDDBUF_6 RE_LU1 
+ RE_RU1 RW_RE_5 RW_RE_6 SAEB_LU1 SAEB_RU1 VDDHD VDDI VSSI WE_LU1 WE_RU1 
+ NET228 WLPYB_6 NET226 WLPY_6 WLP_SAE_5 WLP_SAE_TK_5 WLP_SAE_TK_6 WLP_SAE_6 
+ YL_5[0] YL_LU1[0] YL_LU1[1] YL_RU1[0] YL_RU1[1] YL_6[0] S1AHSF400W40_BK_LCNT_U_SIM
XBK_WLDV_LD_D VDDHD VDDI DEC_X0_2[0] DEC_X0_2[1] DEC_X0_2[2] DEC_X0_2[3] 
+ DEC_X0_2[4] DEC_X0_2[5] DEC_X0_2[6] DEC_X0_2[7] DEC_X0_3[0] DEC_X0_3[1] 
+ DEC_X0_3[2] DEC_X0_3[3] DEC_X0_3[4] DEC_X0_3[5] DEC_X0_3[6] DEC_X0_3[7] 
+ DEC_X1_2[0] DEC_X1_2[1] DEC_X1_2[2] DEC_X1_2[3] DEC_X1_2[4] DEC_X1_2[5] 
+ DEC_X1_2[6] DEC_X1_2[7] DEC_X1_3[0] DEC_X1_3[1] DEC_X1_3[2] DEC_X1_3[3] 
+ DEC_X1_3[4] DEC_X1_3[5] DEC_X1_3[6] DEC_X1_3[7] DEC_X2_2[0] DEC_X2_2[1] 
+ DEC_X2_2[2] DEC_X2_2[3] DEC_X2_3[0] DEC_X2_3[1] DEC_X2_3[2] DEC_X2_3[3] 
+ DEC_X3_2[0] DEC_X3_2[1] DEC_X3_2[2] DEC_X3_2[3] DEC_X3_2[4] DEC_X3_2[5] 
+ DEC_X3_2[6] DEC_X3_2[7] DEC_X3_3[0] DEC_X3_3[1] DEC_X3_3[2] DEC_X3_3[3] 
+ DEC_X3_3[4] DEC_X3_3[5] DEC_X3_3[6] DEC_X3_3[7] DEC_Y_2[0] DEC_Y_2[1] 
+ DEC_Y_2[2] DEC_Y_2[3] DEC_Y_2[4] DEC_Y_2[5] DEC_Y_2[6] DEC_Y_2[7] DEC_Y_3[0] 
+ DEC_Y_3[1] DEC_Y_3[2] DEC_Y_3[3] DEC_Y_3[4] DEC_Y_3[5] DEC_Y_3[6] DEC_Y_3[7] 
+ PD_BUF_2 PD_BUF_3 PD_CVDDBUF_2 PD_CVDDBUF_3 RW_RE_2 RW_RE_3 VDDHD VDDI VSSI 
+ WLP_SAE_2 WLP_SAE_TK_2 WLP_SAE_TK_3 WLP_SAE_3 YL_2[0] YL_3[0] 
+ S1AHSF400W40_BK_WLDV_LD_SIM
XBK_WLDV_LD_U VDDHD VDDI DEC_X0_6[0] DEC_X0_6[1] DEC_X0_6[2] DEC_X0_6[3] 
+ DEC_X0_6[4] DEC_X0_6[5] DEC_X0_6[6] DEC_X0_6[7] DEC_X0_7[0] DEC_X0_7[1] 
+ DEC_X0_7[2] DEC_X0_7[3] DEC_X0_7[4] DEC_X0_7[5] DEC_X0_7[6] DEC_X0_7[7] 
+ DEC_X1_6[0] DEC_X1_6[1] DEC_X1_6[2] DEC_X1_6[3] DEC_X1_6[4] DEC_X1_6[5] 
+ DEC_X1_6[6] DEC_X1_6[7] DEC_X1_7[0] DEC_X1_7[1] DEC_X1_7[2] DEC_X1_7[3] 
+ DEC_X1_7[4] DEC_X1_7[5] DEC_X1_7[6] DEC_X1_7[7] DEC_X2_6[0] DEC_X2_6[1] 
+ DEC_X2_6[2] DEC_X2_6[3] DEC_X2_7[0] DEC_X2_7[1] DEC_X2_7[2] DEC_X2_7[3] 
+ DEC_X3_6[0] DEC_X3_6[1] DEC_X3_6[2] DEC_X3_6[3] DEC_X3_6[4] DEC_X3_6[5] 
+ DEC_X3_6[6] DEC_X3_6[7] DEC_X3_7[0] DEC_X3_7[1] DEC_X3_7[2] DEC_X3_7[3] 
+ DEC_X3_7[4] DEC_X3_7[5] DEC_X3_7[6] DEC_X3_7[7] DEC_Y_6[0] DEC_Y_6[1] 
+ DEC_Y_6[2] DEC_Y_6[3] DEC_Y_6[4] DEC_Y_6[5] DEC_Y_6[6] DEC_Y_6[7] DEC_Y_7[0] 
+ DEC_Y_7[1] DEC_Y_7[2] DEC_Y_7[3] DEC_Y_7[4] DEC_Y_7[5] DEC_Y_7[6] DEC_Y_7[7] 
+ PD_BUF_6 PD_BUF_7 PD_CVDDBUF_6 PD_CVDDBUF_7 RW_RE_6 RW_RE_7 VDDHD VDDI VSSI 
+ WLP_SAE_6 WLP_SAE_TK_6 WLP_SAE_TK_7 WLP_SAE_7 YL_6[0] YL_7[0] 
+ S1AHSF400W40_BK_WLDV_LD_SIM
XTRKPRE PD TRKBL WL_TK VDDHD VDDI VSSI TIEH_BT TIEL S1AHSF400W40_TRKPRE_SIM
XBK_TOP_EDGE VDDHD VDDI VSSI WLP_SAE_8 WLP_SAE_TK_8 S1AHSF400W40_BK_TOP_EDGE_SIM
XARR_LIO_LD_RU BLEQ_DN_RU2 BLEQ_DN_RU3 BLEQ_UP_RU2 BLEQ_UP_RU3 VDDI RE_RU2 
+ RE_RU3 SAEB_RU2 SAEB_RU3 VDDHD VDDI VSSI WE_RU2 WE_RU3 YL_RU2[0] YL_RU2[1] 
+ YL_RU3[0] YL_RU3[1] Y_DN_RU2[0] Y_DN_RU2[1] Y_DN_RU2[2] Y_DN_RU2[3] 
+ Y_DN_RU2[4] Y_DN_RU2[5] Y_DN_RU2[6] Y_DN_RU2[7] Y_DN_RU3[0] Y_DN_RU3[1] 
+ Y_DN_RU3[2] Y_DN_RU3[3] Y_DN_RU3[4] Y_DN_RU3[5] Y_DN_RU3[6] Y_DN_RU3[7] 
+ Y_UP_RU2[0] Y_UP_RU2[1] Y_UP_RU2[2] Y_UP_RU2[3] Y_UP_RU2[4] Y_UP_RU2[5] 
+ Y_UP_RU2[6] Y_UP_RU2[7] Y_UP_RU3[0] Y_UP_RU3[1] Y_UP_RU3[2] Y_UP_RU3[3] 
+ Y_UP_RU3[4] Y_UP_RU3[5] Y_UP_RU3[6] Y_UP_RU3[7] S1AHSF400W40_ARR_LIO_LD_SIM
XARR_LIO_LD_LD BLEQ_DN_LD3 BLEQ_DN_LD2 BLEQ_UP_LD3 BLEQ_UP_LD2 VDDI RE_LD3 
+ RE_LD2 SAEB_LD3 SAEB_LD2 VDDHD VDDI VSSI WE_LD3 WE_LD2 YL_LD3[0] YL_LD3[1] 
+ YL_LD2[0] YL_LD2[1] Y_DN_LD3[0] Y_DN_LD3[1] Y_DN_LD3[2] Y_DN_LD3[3] 
+ Y_DN_LD3[4] Y_DN_LD3[5] Y_DN_LD3[6] Y_DN_LD3[7] Y_DN_LD2[0] Y_DN_LD2[1] 
+ Y_DN_LD2[2] Y_DN_LD2[3] Y_DN_LD2[4] Y_DN_LD2[5] Y_DN_LD2[6] Y_DN_LD2[7] 
+ Y_UP_LD3[0] Y_UP_LD3[1] Y_UP_LD3[2] Y_UP_LD3[3] Y_UP_LD3[4] Y_UP_LD3[5] 
+ Y_UP_LD3[6] Y_UP_LD3[7] Y_UP_LD2[0] Y_UP_LD2[1] Y_UP_LD2[2] Y_UP_LD2[3] 
+ Y_UP_LD2[4] Y_UP_LD2[5] Y_UP_LD2[6] Y_UP_LD2[7] S1AHSF400W40_ARR_LIO_LD_SIM
XARR_LIO_LD_RD BLEQ_DN_RD2 BLEQ_DN_RD3 BLEQ_UP_RD2 BLEQ_UP_RD3 VDDI RE_RD2 
+ RE_RD3 SAEB_RD2 SAEB_RD3 VDDHD VDDI VSSI WE_RD2 WE_RD3 YL_RD2[0] YL_RD2[1] 
+ YL_RD3[0] YL_RD3[1] Y_DN_RD2[0] Y_DN_RD2[1] Y_DN_RD2[2] Y_DN_RD2[3] 
+ Y_DN_RD2[4] Y_DN_RD2[5] Y_DN_RD2[6] Y_DN_RD2[7] Y_DN_RD3[0] Y_DN_RD3[1] 
+ Y_DN_RD3[2] Y_DN_RD3[3] Y_DN_RD3[4] Y_DN_RD3[5] Y_DN_RD3[6] Y_DN_RD3[7] 
+ Y_UP_RD2[0] Y_UP_RD2[1] Y_UP_RD2[2] Y_UP_RD2[3] Y_UP_RD2[4] Y_UP_RD2[5] 
+ Y_UP_RD2[6] Y_UP_RD2[7] Y_UP_RD3[0] Y_UP_RD3[1] Y_UP_RD3[2] Y_UP_RD3[3] 
+ Y_UP_RD3[4] Y_UP_RD3[5] Y_UP_RD3[6] Y_UP_RD3[7] S1AHSF400W40_ARR_LIO_LD_SIM
XARR_LIO_LD_LU BLEQ_DN_LU3 BLEQ_DN_LU2 BLEQ_UP_LU3 BLEQ_UP_LU2 VDDI RE_LU3 
+ RE_LU2 SAEB_LU3 SAEB_LU2 VDDHD VDDI VSSI WE_LU3 WE_LU2 YL_LU3[0] YL_LU3[1] 
+ YL_LU2[0] YL_LU2[1] Y_DN_LU3[0] Y_DN_LU3[1] Y_DN_LU3[2] Y_DN_LU3[3] 
+ Y_DN_LU3[4] Y_DN_LU3[5] Y_DN_LU3[6] Y_DN_LU3[7] Y_DN_LU2[0] Y_DN_LU2[1] 
+ Y_DN_LU2[2] Y_DN_LU2[3] Y_DN_LU2[4] Y_DN_LU2[5] Y_DN_LU2[6] Y_DN_LU2[7] 
+ Y_UP_LU3[0] Y_UP_LU3[1] Y_UP_LU3[2] Y_UP_LU3[3] Y_UP_LU3[4] Y_UP_LU3[5] 
+ Y_UP_LU3[6] Y_UP_LU3[7] Y_UP_LU2[0] Y_UP_LU2[1] Y_UP_LU2[2] Y_UP_LU2[3] 
+ Y_UP_LU2[4] Y_UP_LU2[5] Y_UP_LU2[6] Y_UP_LU2[7] S1AHSF400W40_ARR_LIO_LD_SIM
XARR_LIO_RUL NET1201 NET0410 NET0411[0] NET0411[1] NET0411[2] NET0411[3] 
+ NET0411[4] NET0411[5] NET0411[6] NET0411[7] NET0411[8] NET0411[9] 
+ NET0411[10] NET0411[11] NET0411[12] NET0411[13] NET428 NET0412 NET0413[0] 
+ NET0413[1] NET0413[2] NET0413[3] NET0413[4] NET0413[5] NET0413[6] NET0413[7] 
+ NET0413[8] NET0413[9] NET0413[10] NET0413[11] NET0413[12] NET0413[13] 
+ BLEQ_DN_RU1 BLEQ_DN_RU2 BLEQ_UP_RU1 BLEQ_UP_RU2 NET1185 NET0417 NET0416[0] 
+ NET0416[1] NET0416[2] NET0416[3] NET0416[4] NET0416[5] NET0416[6] NET0416[7] 
+ NET0416[8] NET0416[9] NET0416[10] NET0416[11] NET0416[12] NET0416[13] 
+ NET1157 NET0415 NET0414[0] NET0414[1] NET0414[2] NET0414[3] NET0414[4] 
+ NET0414[5] NET0414[6] NET0414[7] NET0414[8] NET0414[9] NET0414[10] 
+ NET0414[11] NET0414[12] NET0414[13] VDDI NET434 NET433 NET432 NET431 NET430 
+ NET429 NET1237 NET1175 RE_RU1 RE_RU2 SAEB_RU1 SAEB_RU2 VDDHD VDDI VSSI 
+ WE_RU1 WE_RU2 YL_RU1[0] YL_RU1[1] YL_RU2[0] YL_RU2[1] Y_DN_RU1[0] 
+ Y_DN_RU1[1] Y_DN_RU1[2] Y_DN_RU1[3] Y_DN_RU1[4] Y_DN_RU1[5] Y_DN_RU1[6] 
+ Y_DN_RU1[7] Y_DN_RU2[0] Y_DN_RU2[1] Y_DN_RU2[2] Y_DN_RU2[3] Y_DN_RU2[4] 
+ Y_DN_RU2[5] Y_DN_RU2[6] Y_DN_RU2[7] Y_UP_RU1[0] Y_UP_RU1[1] Y_UP_RU1[2] 
+ Y_UP_RU1[3] Y_UP_RU1[4] Y_UP_RU1[5] Y_UP_RU1[6] Y_UP_RU1[7] Y_UP_RU2[0] 
+ Y_UP_RU2[1] Y_UP_RU2[2] Y_UP_RU2[3] Y_UP_RU2[4] Y_UP_RU2[5] Y_UP_RU2[6] 
+ Y_UP_RU2[7] S1AHSF400W40_ARR_LIO_SIM
XARR_LIO_RUR NET1179 NET0450 NET0451[0] NET0451[1] NET0451[2] NET0451[3] 
+ NET0451[4] NET0451[5] NET0451[6] NET0451[7] NET0451[8] NET0451[9] 
+ NET0451[10] NET0451[11] NET0451[12] NET0451[13] NET1167 NET0452 NET0453[0] 
+ NET0453[1] NET0453[2] NET0453[3] NET0453[4] NET0453[5] NET0453[6] NET0453[7] 
+ NET0453[8] NET0453[9] NET0453[10] NET0453[11] NET0453[12] NET0453[13] 
+ BLEQ_DN_RU3 BLEQ_DN_RU4 BLEQ_UP_RU3 BLEQ_UP_RU4 NET1196 NET0457 NET0456[0] 
+ NET0456[1] NET0456[2] NET0456[3] NET0456[4] NET0456[5] NET0456[6] NET0456[7] 
+ NET0456[8] NET0456[9] NET0456[10] NET0456[11] NET0456[12] NET0456[13] 
+ NET1150 NET0455 NET0454[0] NET0454[1] NET0454[2] NET0454[3] NET0454[4] 
+ NET0454[5] NET0454[6] NET0454[7] NET0454[8] NET0454[9] NET0454[10] 
+ NET0454[11] NET0454[12] NET0454[13] VDDI NET1238 NET1219 NET1262 NET1261 
+ NET1126 NET1174 NET1137 NET1254 RE_RU3 RE_RU4 SAEB_RU3 SAEB_RU4 VDDHD VDDI 
+ VSSI WE_RU3 WE_RU4 YL_RU3[0] YL_RU3[1] YL_RU4[0] YL_RU4[1] Y_DN_RU3[0] 
+ Y_DN_RU3[1] Y_DN_RU3[2] Y_DN_RU3[3] Y_DN_RU3[4] Y_DN_RU3[5] Y_DN_RU3[6] 
+ Y_DN_RU3[7] Y_DN_RU4[0] Y_DN_RU4[1] Y_DN_RU4[2] Y_DN_RU4[3] Y_DN_RU4[4] 
+ Y_DN_RU4[5] Y_DN_RU4[6] Y_DN_RU4[7] Y_UP_RU3[0] Y_UP_RU3[1] Y_UP_RU3[2] 
+ Y_UP_RU3[3] Y_UP_RU3[4] Y_UP_RU3[5] Y_UP_RU3[6] Y_UP_RU3[7] Y_UP_RU4[0] 
+ Y_UP_RU4[1] Y_UP_RU4[2] Y_UP_RU4[3] Y_UP_RU4[4] Y_UP_RU4[5] Y_UP_RU4[6] 
+ Y_UP_RU4[7] S1AHSF400W40_ARR_LIO_SIM
XARR_LIO_LDR BLB_LR_3 BLB_DUM_LR_3 NET0491[0] NET0491[1] NET0491[2] NET0491[3] 
+ NET0491[4] NET0491[5] NET0491[6] NET0491[7] NET0491[8] NET0491[9] 
+ NET0491[10] NET0491[11] NET0491[12] NET0491[13] NET1224 NET0492 NET0493[0] 
+ NET0493[1] NET0493[2] NET0493[3] NET0493[4] NET0493[5] NET0493[6] NET0493[7] 
+ NET0493[8] NET0493[9] NET0493[10] NET0493[11] NET0493[12] NET0493[13] 
+ BLEQ_DN_LD2 BLEQ_DN_LD1 BLEQ_UP_LD2 BLEQ_UP_LD1 BL_LR_3 BL_DUM_LR_3 
+ NET0496[0] NET0496[1] NET0496[2] NET0496[3] NET0496[4] NET0496[5] NET0496[6] 
+ NET0496[7] NET0496[8] NET0496[9] NET0496[10] NET0496[11] NET0496[12] 
+ NET0496[13] NET1205 NET0495 NET0494[0] NET0494[1] NET0494[2] NET0494[3] 
+ NET0494[4] NET0494[5] NET0494[6] NET0494[7] NET0494[8] NET0494[9] 
+ NET0494[10] NET0494[11] NET0494[12] NET0494[13] VDDI GBLB_LR_3 GBLB_LR_4 
+ GBL_LR_3 GBL_LR_4 GWB_LR_3 GWB_LR_4 GW_LR_3 GW_LR_4 RE_LD2 RE_LD1 SAEB_LD2 
+ SAEB_LD1 VDDHD VDDI VSSI WE_LD2 WE_LD1 YL_LD2[0] YL_LD2[1] YL_LD1[0] 
+ YL_LD1[1] Y_DN_LD2[0] Y_DN_LD2[1] Y_DN_LD2[2] Y_DN_LD2[3] Y_DN_LD2[4] 
+ Y_DN_LD2[5] Y_DN_LD2[6] Y_DN_LD2[7] Y_DN_LD1[0] Y_DN_LD1[1] Y_DN_LD1[2] 
+ Y_DN_LD1[3] Y_DN_LD1[4] Y_DN_LD1[5] Y_DN_LD1[6] Y_DN_LD1[7] Y_UP_LD2[0] 
+ Y_UP_LD2[1] Y_UP_LD2[2] Y_UP_LD2[3] Y_UP_LD2[4] Y_UP_LD2[5] Y_UP_LD2[6] 
+ Y_UP_LD2[7] Y_UP_LD1[0] Y_UP_LD1[1] Y_UP_LD1[2] Y_UP_LD1[3] Y_UP_LD1[4] 
+ Y_UP_LD1[5] Y_UP_LD1[6] Y_UP_LD1[7] S1AHSF400W40_ARR_LIO_SIM
XARR_LIO_RDR NET527 NET0530 NET0531[0] NET0531[1] NET0531[2] NET0531[3] 
+ NET0531[4] NET0531[5] NET0531[6] NET0531[7] NET0531[8] NET0531[9] 
+ NET0531[10] NET0531[11] NET0531[12] NET0531[13] NET536 NET0532 NET0533[0] 
+ NET0533[1] NET0533[2] NET0533[3] NET0533[4] NET0533[5] NET0533[6] NET0533[7] 
+ NET0533[8] NET0533[9] NET0533[10] NET0533[11] NET0533[12] NET0533[13] 
+ BLEQ_DN_RD3 BLEQ_DN_RD4 BLEQ_UP_RD3 BLEQ_UP_RD4 NET535 NET0537 NET0536[0] 
+ NET0536[1] NET0536[2] NET0536[3] NET0536[4] NET0536[5] NET0536[6] NET0536[7] 
+ NET0536[8] NET0536[9] NET0536[10] NET0536[11] NET0536[12] NET0536[13] NET531 
+ NET0535 NET0534[0] NET0534[1] NET0534[2] NET0534[3] NET0534[4] NET0534[5] 
+ NET0534[6] NET0534[7] NET0534[8] NET0534[9] NET0534[10] NET0534[11] 
+ NET0534[12] NET0534[13] VDDI NET542 NET541 NET540 NET539 NET538 NET537 
+ NET534 NET533 RE_RD3 RE_RD4 SAEB_RD3 SAEB_RD4 VDDHD VDDI VSSI WE_RD3 WE_RD4 
+ YL_RD3[0] YL_RD3[1] YL_RD4[0] YL_RD4[1] Y_DN_RD3[0] Y_DN_RD3[1] Y_DN_RD3[2] 
+ Y_DN_RD3[3] Y_DN_RD3[4] Y_DN_RD3[5] Y_DN_RD3[6] Y_DN_RD3[7] Y_DN_RD4[0] 
+ Y_DN_RD4[1] Y_DN_RD4[2] Y_DN_RD4[3] Y_DN_RD4[4] Y_DN_RD4[5] Y_DN_RD4[6] 
+ Y_DN_RD4[7] Y_UP_RD3[0] Y_UP_RD3[1] Y_UP_RD3[2] Y_UP_RD3[3] Y_UP_RD3[4] 
+ Y_UP_RD3[5] Y_UP_RD3[6] Y_UP_RD3[7] Y_UP_RD4[0] Y_UP_RD4[1] Y_UP_RD4[2] 
+ Y_UP_RD4[3] Y_UP_RD4[4] Y_UP_RD4[5] Y_UP_RD4[6] Y_UP_RD4[7] S1AHSF400W40_ARR_LIO_SIM
XARR_LIO_RDL NET1162 NET0570 NET0571[0] NET0571[1] NET0571[2] NET0571[3] 
+ NET0571[4] NET0571[5] NET0571[6] NET0571[7] NET0571[8] NET0571[9] 
+ NET0571[10] NET0571[11] NET0571[12] NET0571[13] NET1135 NET0572 NET0573[0] 
+ NET0573[1] NET0573[2] NET0573[3] NET0573[4] NET0573[5] NET0573[6] NET0573[7] 
+ NET0573[8] NET0573[9] NET0573[10] NET0573[11] NET0573[12] NET0573[13] 
+ BLEQ_DN_RD1 BLEQ_DN_RD2 BLEQ_UP_RD1 BLEQ_UP_RD2 NET1249 NET0577 NET0576[0] 
+ NET0576[1] NET0576[2] NET0576[3] NET0576[4] NET0576[5] NET0576[6] NET0576[7] 
+ NET0576[8] NET0576[9] NET0576[10] NET0576[11] NET0576[12] NET0576[13] 
+ NET1156 NET0575 NET0574[0] NET0574[1] NET0574[2] NET0574[3] NET0574[4] 
+ NET0574[5] NET0574[6] NET0574[7] NET0574[8] NET0574[9] NET0574[10] 
+ NET0574[11] NET0574[12] NET0574[13] VDDI NET1255 NET1266 NET1190 NET1264 
+ NET1231 NET1270 NET1163 NET1109 RE_RD1 RE_RD2 SAEB_RD1 SAEB_RD2 VDDHD VDDI 
+ VSSI WE_RD1 WE_RD2 YL_RD1[0] YL_RD1[1] YL_RD2[0] YL_RD2[1] Y_DN_RD1[0] 
+ Y_DN_RD1[1] Y_DN_RD1[2] Y_DN_RD1[3] Y_DN_RD1[4] Y_DN_RD1[5] Y_DN_RD1[6] 
+ Y_DN_RD1[7] Y_DN_RD2[0] Y_DN_RD2[1] Y_DN_RD2[2] Y_DN_RD2[3] Y_DN_RD2[4] 
+ Y_DN_RD2[5] Y_DN_RD2[6] Y_DN_RD2[7] Y_UP_RD1[0] Y_UP_RD1[1] Y_UP_RD1[2] 
+ Y_UP_RD1[3] Y_UP_RD1[4] Y_UP_RD1[5] Y_UP_RD1[6] Y_UP_RD1[7] Y_UP_RD2[0] 
+ Y_UP_RD2[1] Y_UP_RD2[2] Y_UP_RD2[3] Y_UP_RD2[4] Y_UP_RD2[5] Y_UP_RD2[6] 
+ Y_UP_RD2[7] S1AHSF400W40_ARR_LIO_SIM
XARR_LIO_LDL BLB_LL_3 BLB_DUM_LL3 NET0611[0] NET0611[1] NET0611[2] NET0611[3] 
+ NET0611[4] NET0611[5] NET0611[6] NET0611[7] NET0611[8] NET0611[9] 
+ NET0611[10] NET0611[11] NET0611[12] NET0611[13] NET1233 NET0612 NET0613[0] 
+ NET0613[1] NET0613[2] NET0613[3] NET0613[4] NET0613[5] NET0613[6] NET0613[7] 
+ NET0613[8] NET0613[9] NET0613[10] NET0613[11] NET0613[12] NET0613[13] 
+ BLEQ_DN_LD4 BLEQ_DN_LD3 BLEQ_UP_LD4 BLEQ_UP_LD3 BL_LL_3 BL_DUM_LL_3 
+ NET0616[0] NET0616[1] NET0616[2] NET0616[3] NET0616[4] NET0616[5] NET0616[6] 
+ NET0616[7] NET0616[8] NET0616[9] NET0616[10] NET0616[11] NET0616[12] 
+ NET0616[13] NET1227 NET0615 NET0614[0] NET0614[1] NET0614[2] NET0614[3] 
+ NET0614[4] NET0614[5] NET0614[6] NET0614[7] NET0614[8] NET0614[9] 
+ NET0614[10] NET0614[11] NET0614[12] NET0614[13] VDDI GBLB_LL_3 GBLB_LL_4 
+ GBL_LL_3 GBL_LL_4 GWB_LL_3 GWB_LL_4 GW_LL_3 GW_LL_4 RE_LD4 RE_LD3 SAEB_LD4 
+ SAEB_LD3 VDDHD VDDI VSSI WE_LD4 WE_LD3 YL_LD4[0] YL_LD4[1] YL_LD3[0] 
+ YL_LD3[1] Y_DN_LD4[0] Y_DN_LD4[1] Y_DN_LD4[2] Y_DN_LD4[3] Y_DN_LD4[4] 
+ Y_DN_LD4[5] Y_DN_LD4[6] Y_DN_LD4[7] Y_DN_LD3[0] Y_DN_LD3[1] Y_DN_LD3[2] 
+ Y_DN_LD3[3] Y_DN_LD3[4] Y_DN_LD3[5] Y_DN_LD3[6] Y_DN_LD3[7] Y_UP_LD4[0] 
+ Y_UP_LD4[1] Y_UP_LD4[2] Y_UP_LD4[3] Y_UP_LD4[4] Y_UP_LD4[5] Y_UP_LD4[6] 
+ Y_UP_LD4[7] Y_UP_LD3[0] Y_UP_LD3[1] Y_UP_LD3[2] Y_UP_LD3[3] Y_UP_LD3[4] 
+ Y_UP_LD3[5] Y_UP_LD3[6] Y_UP_LD3[7] S1AHSF400W40_ARR_LIO_SIM
XARR_LIO_LUL NET1124 NET0650 NET0651[0] NET0651[1] NET0651[2] NET0651[3] 
+ NET0651[4] NET0651[5] NET0651[6] NET0651[7] NET0651[8] NET0651[9] 
+ NET0651[10] NET0651[11] NET0651[12] NET0651[13] BLB_LL_6 BLB_DUM_LL_6 
+ NET0653[0] NET0653[1] NET0653[2] NET0653[3] NET0653[4] NET0653[5] NET0653[6] 
+ NET0653[7] NET0653[8] NET0653[9] NET0653[10] NET0653[11] NET0653[12] 
+ NET0653[13] BLEQ_DN_LU4 BLEQ_DN_LU3 BLEQ_UP_LU4 BLEQ_UP_LU3 NET1123 NET0657 
+ NET0656[0] NET0656[1] NET0656[2] NET0656[3] NET0656[4] NET0656[5] NET0656[6] 
+ NET0656[7] NET0656[8] NET0656[9] NET0656[10] NET0656[11] NET0656[12] 
+ NET0656[13] BL_LL_6 BL_DUM_LL_6 NET0654[0] NET0654[1] NET0654[2] NET0654[3] 
+ NET0654[4] NET0654[5] NET0654[6] NET0654[7] NET0654[8] NET0654[9] 
+ NET0654[10] NET0654[11] NET0654[12] NET0654[13] VDDI GBLB_LL_5 GBLB_LL_6 
+ GBL_LL_5 GBL_LL_6 GWB_LL_5 GWB_LL_6 GW_LL_5 GW_LL_6 RE_LU4 RE_LU3 SAEB_LU4 
+ SAEB_LU3 VDDHD VDDI VSSI WE_LU4 WE_LU3 YL_LU4[0] YL_LU4[1] YL_LU3[0] 
+ YL_LU3[1] Y_DN_LU4[0] Y_DN_LU4[1] Y_DN_LU4[2] Y_DN_LU4[3] Y_DN_LU4[4] 
+ Y_DN_LU4[5] Y_DN_LU4[6] Y_DN_LU4[7] Y_DN_LU3[0] Y_DN_LU3[1] Y_DN_LU3[2] 
+ Y_DN_LU3[3] Y_DN_LU3[4] Y_DN_LU3[5] Y_DN_LU3[6] Y_DN_LU3[7] Y_UP_LU4[0] 
+ Y_UP_LU4[1] Y_UP_LU4[2] Y_UP_LU4[3] Y_UP_LU4[4] Y_UP_LU4[5] Y_UP_LU4[6] 
+ Y_UP_LU4[7] Y_UP_LU3[0] Y_UP_LU3[1] Y_UP_LU3[2] Y_UP_LU3[3] Y_UP_LU3[4] 
+ Y_UP_LU3[5] Y_UP_LU3[6] Y_UP_LU3[7] S1AHSF400W40_ARR_LIO_SIM
XARR_LIO_LUR NET1191 NET0690 NET0691[0] NET0691[1] NET0691[2] NET0691[3] 
+ NET0691[4] NET0691[5] NET0691[6] NET0691[7] NET0691[8] NET0691[9] 
+ NET0691[10] NET0691[11] NET0691[12] NET0691[13] BLB_LR_6 BLB_DUM_LR_6 
+ NET0693[0] NET0693[1] NET0693[2] NET0693[3] NET0693[4] NET0693[5] NET0693[6] 
+ NET0693[7] NET0693[8] NET0693[9] NET0693[10] NET0693[11] NET0693[12] 
+ NET0693[13] BLEQ_DN_LU2 BLEQ_DN_LU1 BLEQ_UP_LU2 BLEQ_UP_LU1 NET1206 NET0697 
+ NET0696[0] NET0696[1] NET0696[2] NET0696[3] NET0696[4] NET0696[5] NET0696[6] 
+ NET0696[7] NET0696[8] NET0696[9] NET0696[10] NET0696[11] NET0696[12] 
+ NET0696[13] BL_LR_6 BL_DUM_LR_6 NET0694[0] NET0694[1] NET0694[2] NET0694[3] 
+ NET0694[4] NET0694[5] NET0694[6] NET0694[7] NET0694[8] NET0694[9] 
+ NET0694[10] NET0694[11] NET0694[12] NET0694[13] VDDI GBLB_LR_5 GBLB_LR_6 
+ GBL_LR_5 GBL_LR_6 GWB_LR_5 GWB_LR_6 GW_LR_5 GW_LR_6 RE_LU2 RE_LU1 SAEB_LU2 
+ SAEB_LU1 VDDHD VDDI VSSI WE_LU2 WE_LU1 YL_LU2[0] YL_LU2[1] YL_LU1[0] 
+ YL_LU1[1] Y_DN_LU2[0] Y_DN_LU2[1] Y_DN_LU2[2] Y_DN_LU2[3] Y_DN_LU2[4] 
+ Y_DN_LU2[5] Y_DN_LU2[6] Y_DN_LU2[7] Y_DN_LU1[0] Y_DN_LU1[1] Y_DN_LU1[2] 
+ Y_DN_LU1[3] Y_DN_LU1[4] Y_DN_LU1[5] Y_DN_LU1[6] Y_DN_LU1[7] Y_UP_LU2[0] 
+ Y_UP_LU2[1] Y_UP_LU2[2] Y_UP_LU2[3] Y_UP_LU2[4] Y_UP_LU2[5] Y_UP_LU2[6] 
+ Y_UP_LU2[7] Y_UP_LU1[0] Y_UP_LU1[1] Y_UP_LU1[2] Y_UP_LU1[3] Y_UP_LU1[4] 
+ Y_UP_LU1[5] Y_UP_LU1[6] Y_UP_LU1[7] S1AHSF400W40_ARR_LIO_SIM
XARR_SEG_LD_LR VDDI GBLB_LR_4 GBLB_LR_5 GBL_LR_4 GBL_LR_5 GWB_LR_4 GWB_LR_5 
+ GW_LR_4 GW_LR_5 VDDHD VDDI VSSI S1AHSF400W40_ARR_SEG_LD_SIM
XARR_SEG_LD_LL VDDI GBLB_LL_4 GBLB_LL_5 GBL_LL_4 GBL_LL_5 GWB_LL_4 GWB_LL_5 
+ GW_LL_4 GW_LL_5 VDDHD VDDI VSSI S1AHSF400W40_ARR_SEG_LD_SIM
XARR_MCB_RUR NET01237 NET01244 NET01242 NET01235 VDDI NET01231 NET01240 
+ NET01238 NET01233 VDDHD VDDI VSSI WL_RU3[0] WL_RU3[1] WL_RU4[0] WL_RU4[1] 
+ S1AHSF400W40_ARR_MCB_SIM
XARR_MCB_RUL NET01254 NET01257 NET01255 NET01256 VDDI NET01260 NET01261 
+ NET01259 NET01258 VDDHD VDDI VSSI WL_RU1[0] WL_RU1[1] WL_RU2[0] WL_RU2[1] 
+ S1AHSF400W40_ARR_MCB_SIM
XARR_MCB_LUR BL_LR_7 BL_DUM_LR_7 BLB_LR_7 BLB_DUM_LR_7 VDDI GBL_LR_78 
+ GBLB_LR_78 GW_LR_78 GWB_LR_78 VDDHD VDDI VSSI WL_LU2[0] WL_LU2[1] WL_LU1[0] 
+ WL_LU1[1] S1AHSF400W40_ARR_MCB_SIM
XARR_MCB_LDL BL_LL_2 BL_DUM_LL_2 BLB_LL_2 BLB_DUM_LL_2 VDDI GBL_LL_12 
+ GBLB_LL_12 GW_LL_12 GWB_LL_12 VDDHD VDDI VSSI WL_LD4[0] WL_LD4[1] WL_LD3[0] 
+ WL_LD3[1] S1AHSF400W40_ARR_MCB_SIM
XARR_MCB_RDR NET01216 NET01225 NET01223 NET01214 VDDI NET01218 NET01219 
+ NET01221 NET01226 VDDHD VDDI VSSI WL_RD3[0] WL_RD3[1] WL_RD4[0] WL_RD4[1] 
+ S1AHSF400W40_ARR_MCB_SIM
XARR_MCB_LDR BL_LR_2 BL_DUM_LR_2 BLB_LR_2 BLB_DUM_LR_2 VDDI GBL_LR_12 
+ GBLB_LR_12 GW_LR_12 GWB_LR_12 VDDHD VDDI VSSI WL_LD2[0] WL_LD2[1] WL_LD1[0] 
+ WL_LD1[1] S1AHSF400W40_ARR_MCB_SIM
XARR_MCB_LUL BL_LL_7 BL_DUM_LL_7 BLB_LL_7 BLB_DUM_LL_7 VDDI GBL_LL_78 
+ GBLB_LL_78 GW_LL_78 GWB_LL_78 VDDHD VDDI VSSI WL_LU4[0] WL_LU4[1] WL_LU3[0] 
+ WL_LU3[1] S1AHSF400W40_ARR_MCB_SIM
XARR_MCB_RDL NET01211 NET01212 NET01210 NET01213 VDDI NET01199 NET01198 
+ NET01206 NET01207 VDDHD VDDI VSSI WL_RD1[0] WL_RD1[1] WL_RD2[0] WL_RD2[1] 
+ S1AHSF400W40_ARR_MCB_SIM
XBK_SEG_LD VDDHD VDDI DEC_X0_4[0] DEC_X0_4[1] DEC_X0_4[2] DEC_X0_4[3] 
+ DEC_X0_4[4] DEC_X0_4[5] DEC_X0_4[6] DEC_X0_4[7] DEC_X0_5[0] DEC_X0_5[1] 
+ DEC_X0_5[2] DEC_X0_5[3] DEC_X0_5[4] DEC_X0_5[5] DEC_X0_5[6] DEC_X0_5[7] 
+ DEC_X1_4[0] DEC_X1_4[1] DEC_X1_4[2] DEC_X1_4[3] DEC_X1_4[4] DEC_X1_4[5] 
+ DEC_X1_4[6] DEC_X1_4[7] DEC_X1_5[0] DEC_X1_5[1] DEC_X1_5[2] DEC_X1_5[3] 
+ DEC_X1_5[4] DEC_X1_5[5] DEC_X1_5[6] DEC_X1_5[7] DEC_X2_4[0] DEC_X2_4[1] 
+ DEC_X2_4[2] DEC_X2_4[3] DEC_X2_5[0] DEC_X2_5[1] DEC_X2_5[2] DEC_X2_5[3] 
+ DEC_X3_4[0] DEC_X3_4[1] DEC_X3_4[2] DEC_X3_4[3] DEC_X3_4[4] DEC_X3_4[5] 
+ DEC_X3_4[6] DEC_X3_4[7] DEC_X3_5[0] DEC_X3_5[1] DEC_X3_5[2] DEC_X3_5[3] 
+ DEC_X3_5[4] DEC_X3_5[5] DEC_X3_5[6] DEC_X3_5[7] DEC_Y_4[0] DEC_Y_4[1] 
+ DEC_Y_4[2] DEC_Y_4[3] DEC_Y_4[4] DEC_Y_4[5] DEC_Y_4[6] DEC_Y_4[7] DEC_Y_5[0] 
+ DEC_Y_5[1] DEC_Y_5[2] DEC_Y_5[3] DEC_Y_5[4] DEC_Y_5[5] DEC_Y_5[6] DEC_Y_5[7] 
+ PD_BUF_4 PD_BUF_5 PD_CVDDBUF_4 PD_CVDDBUF_5 RW_RE_4 RW_RE_5 VDDHD VDDI VSSI 
+ WLP_SAE_4 WLP_SAE_TK_4 WLP_SAE_TK_5 WLP_SAE_5 YL_4[0] YL_5[0] S1AHSF400W40_BK_SEG_LD_SIM
XARR_WLLD_LU VDDI VDDHD VDDI VSSI WL_LU3[0] WL_LU3[1] WL_LU2[0] WL_LU2[1] 
+ S1AHSF400W40_ARR_WLLD_SIM
XARR_WLLD_RU VDDI VDDHD VDDI VSSI WL_RU2[0] WL_RU2[1] WL_RU3[0] WL_RU3[1] 
+ S1AHSF400W40_ARR_WLLD_SIM
XARR_WLLD_LD VDDI VDDHD VDDI VSSI WL_LD3[0] WL_LD3[1] WL_LD2[0] WL_LD2[1] 
+ S1AHSF400W40_ARR_WLLD_SIM
XARR_WLLD_RD VDDI VDDHD VDDI VSSI WL_RD2[0] WL_RD2[1] WL_RD3[0] WL_RD3[1] 
+ S1AHSF400W40_ARR_WLLD_SIM
XARR_BLLD_LUL BLB_LL_6 BLB_DUM_LL_6 BLB_LL_7 BLB_DUM_LL_7 BL_LL_6 BL_DUM_LL_6 
+ BL_LL_7 BL_DUM_LL_7 VDDI GBLB_LL_6 GBLB_LL_78 GBL_LL_6 GBL_LL_78 GWB_LL_6 
+ GWB_LL_78 GW_LL_6 GW_LL_78 VDDHD VDDI VSSI S1AHSF400W40_ARR_BLLD_SIM
XARRLBLLD_LDL BLB_LL_2 BLB_DUM_LL_2 BLB_LL_3 BLB_DUM_LL3 BL_LL_2 BL_DUM_LL_2 
+ BL_LL_3 BL_DUM_LL_3 VDDI GBLB_LL_12 GBLB_LL_3 GBL_LL_12 GBL_LL_3 GWB_LL_12 
+ GWB_LL_3 GW_LL_12 GW_LL_3 VDDHD VDDI VSSI S1AHSF400W40_ARR_BLLD_SIM
XARR_BLLD_LDR BLB_LR_2 BLB_DUM_LR_2 BLB_LR_3 BLB_DUM_LR_3 BL_LR_2 BL_DUM_LR_2 
+ BL_LR_3 BL_DUM_LR_3 VDDI GBLB_LR_12 GBLB_LR_3 GBL_LR_12 GBL_LR_3 GWB_LR_12 
+ GWB_LR_3 GW_LR_12 GW_LR_3 VDDHD VDDI VSSI S1AHSF400W40_ARR_BLLD_SIM
XARR_BLLD_LUR BLB_LR_6 BLB_DUM_LR_6 BLB_LR_7 BLB_DUM_LR_7 BL_LR_6 BL_DUM_LR_6 
+ BL_LR_7 BL_DUM_LR_7 VDDI GBLB_LR_6 GBLB_LR_78 GBL_LR_6 GBL_LR_78 GWB_LR_6 
+ GWB_LR_78 GW_LR_6 GW_LR_78 VDDHD VDDI VSSI S1AHSF400W40_ARR_BLLD_SIM
XTKBL TRKBL BL_TK_TP VDDHD PD VDDHD VDDI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI 
+ VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI VSSI WL_TK_ACT[0] 
+ WL_TK_ACT[1] WL_TK_ACT[2] WL_TK_ACT[3] WL_TK_ACT[4] WL_TK_ACT[5] 
+ WL_TK_ACT[6] WL_TK_ACT[7] WL_TK_ACT[8] WL_TK_ACT[9] WL_TK_ACT[10] 
+ WL_TK_ACT[11] WL_TK_ACT[12] WL_TK_ACT[13] WL_TK_ACT[14] WL_TK_ACT[15] 
+ WL_TK_ACT[16] WL_TK_ACT[17] WL_TK_ACT[18] WL_TK_ACT[19] WL_TK_ACT[20] 
+ WL_TK_ACT[21] WL_TK_ACT[22] WL_TK_ACT[23] WL_TK_ACT[24] WL_TK_ACT[25] 
+ WL_TK_ACT[26] WL_TK_ACT[27] WL_TK_ACT[28] WL_TK_ACT[29] WL_TK_ACT[30] 
+ WL_TK_ACT[31] WL_TK_ACT[32] WL_TK_ACT[33] WL_TK_ACT[34] WL_TK_ACT[35] 
+ WL_TK_ACT[36] WL_TK_ACT[37] WL_TK_ACT[38] WL_TK_ACT[39] WL_TK_ACT[40] 
+ WL_TK_ACT[41] WL_TK_ACT[42] WL_TK_ACT[43] WL_TK_ACT[44] WL_TK_ACT[45] 
+ WL_TK_ACT[46] WL_TK_ACT[47] WL_TK_ACT[48] WL_TK_ACT[49] WL_TK_ACT[50] 
+ WL_TK_ACT[51] WL_TK_ACT[52] WL_TK_ACT[53] WL_TK_ACT[54] WL_TK_ACT[55] 
+ WL_TK_ACT[56] WL_TK_ACT[57] WL_TK_ACT[58] WL_TK_ACT[59] WL_TK_ACT[60] 
+ WL_TK_ACT[61] WL_TK_ACT[62] WL_TK_ACT[63] WL_TK_ACT[64] WL_TK_ACT[65] 
+ WL_TK_ACT[66] WL_TK_ACT[67] WL_TK_ACT[68] WL_TK_ACT[69] WL_TK_ACT[70] 
+ WL_TK_ACT[71] WL_TK_ACT[72] WL_TK_ACT[73] WL_TK_ACT[74] WL_TK_ACT[75] 
+ WL_TK_ACT[76] WL_TK_ACT[77] WL_TK_ACT[78] WL_TK_ACT[79] WL_TK_ACT[80] 
+ WL_TK_ACT[81] WL_TK_ACT[82] WL_TK_ACT[83] WL_TK_ACT[84] WL_TK_ACT[85] 
+ WL_TK_ACT[86] WL_TK_ACT[87] WL_TK_ACT[88] WL_TK_ACT[89] WL_TK_ACT[90] 
+ WL_TK_ACT[91] WL_TK_ACT[92] WL_TK_ACT[93] WL_TK_ACT[94] WL_TK_ACT[95] 
+ WL_TK_ACT[96] WL_TK_ACT[97] WL_TK_ACT[98] WL_TK_ACT[99] WL_TK_ACT[100] 
+ WL_TK_ACT[101] WL_TK_ACT[102] WL_TK_ACT[103] WL_TK_ACT[104] WL_TK_ACT[105] 
+ WL_TK_ACT[106] WL_TK_ACT[107] WL_TK_ACT[108] WL_TK_ACT[109] WL_TK_ACT[110] 
+ WL_TK_ACT[111] WL_TK_ACT[112] WL_TK_ACT[113] WL_TK_ACT[114] WL_TK_ACT[115] 
+ WL_TK_ACT[116] WL_TK_ACT[117] WL_TK_ACT[118] WL_TK_ACT[119] WL_TK_ACT[120] 
+ WL_TK_ACT[121] WL_TK_ACT[122] WL_TK_ACT[123] WL_TK_ACT[124] WL_TK_ACT[125] 
+ WL_TK_ACT[126] WL_TK_ACT[127] WL_TK_ACT[128] WL_TK_ACT[129] WL_TK_ACT[130] 
+ WL_TK_ACT[131] WL_TK_ACT[132] WL_TK_ACT[133] WL_TK_ACT[134] WL_TK_ACT[135] 
+ WL_TK_ACT[136] WL_TK_ACT[137] WL_TK_ACT[138] WL_TK_ACT[139] WL_TK_ACT[140] 
+ WL_TK_ACT[141] WL_TK_ACT[142] WL_TK_ACT[143] WL_TK_ACT[144] WL_TK_ACT[145] 
+ WL_TK_ACT[146] WL_TK_ACT[147] WL_TK_ACT[148] WL_TK_ACT[149] WL_TK_ACT[150] 
+ WL_TK_ACT[151] WL_TK_ACT[152] WL_TK_ACT[153] WL_TK_ACT[154] WL_TK_ACT[155] 
+ WL_TK_ACT[156] WL_TK_ACT[157] WL_TK_ACT[158] WL_TK_ACT[159] WL_TK_ACT[160] 
+ WL_TK_ACT[161] WL_TK_ACT[162] WL_TK_ACT[163] WL_TK_ACT[164] WL_TK_ACT[165] 
+ WL_TK_ACT[166] WL_TK_ACT[167] WL_TK_ACT[168] WL_TK_ACT[169] WL_TK_ACT[170] 
+ WL_TK_ACT[171] WL_TK_ACT[172] WL_TK_ACT[173] WL_TK_ACT[174] WL_TK_ACT[175] 
+ WL_TK_ACT[176] WL_TK_ACT[177] WL_TK_ACT[178] WL_TK_ACT[179] WL_TK_ACT[180] 
+ WL_TK_ACT[181] WL_TK_ACT[182] WL_TK_ACT[183] WL_TK_ACT[184] WL_TK_ACT[185] 
+ WL_TK_ACT[186] WL_TK_ACT[187] WL_TK_ACT[188] WL_TK_ACT[189] WL_TK_ACT[190] 
+ WL_TK_ACT[191] WL_TK_ACT[192] WL_TK_ACT[193] WL_TK_ACT[194] WL_TK_ACT[195] 
+ WL_TK_ACT[196] WL_TK_ACT[197] WL_TK_ACT[198] WL_TK_ACT[199] WL_TK_ACT[200] 
+ WL_TK_ACT[201] WL_TK_ACT[202] WL_TK_ACT[203] WL_TK_ACT[204] WL_TK_ACT[205] 
+ WL_TK_ACT[206] WL_TK_ACT[207] WL_TK_ACT[208] WL_TK_ACT[209] WL_TK_ACT[210] 
+ WL_TK_ACT[211] WL_TK_ACT[212] WL_TK_ACT[213] WL_TK_ACT[214] WL_TK_ACT[215] 
+ WL_TK_ACT[216] WL_TK_ACT[217] WL_TK_ACT[218] WL_TK_ACT[219] WL_TK_ACT[220] 
+ WL_TK_ACT[221] WL_TK_ACT[222] WL_TK_ACT[223] WL_TK_ACT[224] WL_TK_ACT[225] 
+ WL_TK_ACT[226] WL_TK_ACT[227] WL_TK_ACT[228] WL_TK_ACT[229] WL_TK_ACT[230] 
+ WL_TK_ACT[231] WL_TK_ACT[232] WL_TK_ACT[233] WL_TK_ACT[234] WL_TK_ACT[235] 
+ WL_TK_ACT[236] WL_TK_ACT[237] WL_TK_ACT[238] WL_TK_ACT[239] WL_TK_ACT[240] 
+ WL_TK_ACT[241] WL_TK_ACT[242] WL_TK_ACT[243] WL_TK_ACT[244] WL_TK_ACT[245] 
+ WL_TK_ACT[246] WL_TK_ACT[247] WL_TK_ACT[248] WL_TK_ACT[249] WL_TK_ACT[250] 
+ WL_TK_ACT[251] WL_TK_ACT[252] WL_TK_ACT[253] WL_TK_ACT[254] WL_TK_ACT[255] 
+ WL_TK_ACT[256] WL_TK_ACT[257] WL_TK_ACT[258] WL_TK_ACT[259] WL_TK_ACT[260] 
+ WL_TK_ACT[261] WL_TK_ACT[262] WL_TK_ACT[263] WL_TK_ACT[264] WL_TK_ACT[265] 
+ WL_TK_ACT[266] WL_TK_ACT[267] WL_TK_ACT[268] WL_TK_ACT[269] WL_TK_ACT[270] 
+ WL_TK_ACT[271] WL_TK_ACT[272] WL_TK_ACT[273] WL_TK_ACT[274] WL_TK_ACT[275] 
+ WL_TK_ACT[276] WL_TK_ACT[277] WL_TK_ACT[278] WL_TK_ACT[279] WL_TK_ACT[280] 
+ WL_TK_ACT[281] WL_TK_ACT[282] WL_TK_ACT[283] WL_TK_ACT[284] WL_TK_ACT[285] 
+ WL_TK_ACT[286] WL_TK_ACT[287] WL_TK_ACT[288] WL_TK_ACT[289] WL_TK_ACT[290] 
+ WL_TK_ACT[291] WL_TK_ACT[292] WL_TK_ACT[293] WL_TK_ACT[294] WL_TK_ACT[295] 
+ WL_TK_ACT[296] WL_TK_ACT[297] WL_TK_ACT[298] WL_TK_ACT[299] WL_TK_ACT[300] 
+ WL_TK_ACT[301] WL_TK_ACT[302] WL_TK_ACT[303] WL_TK_ACT[304] WL_TK_ACT[305] 
+ WL_TK_ACT[306] WL_TK_ACT[307] WL_TK_ACT[308] WL_TK_ACT[309] WL_TK_ACT[310] 
+ WL_TK_ACT[311] WL_TK_ACT[312] WL_TK_ACT[313] WL_TK_ACT[314] WL_TK_ACT[315] 
+ WL_TK_ACT[316] WL_TK_ACT[317] WL_TK_ACT[318] WL_TK_ACT[319] WL_TK_ACT[320] 
+ WL_TK_ACT[321] WL_TK_ACT[322] WL_TK_ACT[323] WL_TK_ACT[324] WL_TK_ACT[325] 
+ WL_TK_ACT[326] WL_TK_ACT[327] WL_TK_ACT[328] WL_TK_ACT[329] WL_TK_ACT[330] 
+ WL_TK_ACT[331] WL_TK_ACT[332] WL_TK_ACT[333] WL_TK_ACT[334] WL_TK_ACT[335] 
+ WL_TK_ACT[336] WL_TK_ACT[337] WL_TK_ACT[338] WL_TK_ACT[339] WL_TK_ACT[340] 
+ WL_TK_ACT[341] WL_TK_ACT[342] WL_TK_ACT[343] WL_TK_ACT[344] WL_TK_ACT[345] 
+ WL_TK_ACT[346] WL_TK_ACT[347] WL_TK_ACT[348] WL_TK_ACT[349] WL_TK_ACT[350] 
+ WL_TK_ACT[351] WL_TK_ACT[352] WL_TK_ACT[353] WL_TK_ACT[354] WL_TK_ACT[355] 
+ WL_TK_ACT[356] WL_TK_ACT[357] WL_TK_ACT[358] WL_TK_ACT[359] WL_TK_ACT[360] 
+ WL_TK_ACT[361] WL_TK_ACT[362] WL_TK_ACT[363] WL_TK_ACT[364] WL_TK_ACT[365] 
+ WL_TK_ACT[366] WL_TK_ACT[367] WL_TK_ACT[368] WL_TK_ACT[369] WL_TK_ACT[370] 
+ WL_TK_ACT[371] WL_TK_ACT[372] WL_TK_ACT[373] WL_TK_ACT[374] WL_TK_ACT[375] 
+ WL_TK_ACT[376] WL_TK_ACT[377] WL_TK_ACT[378] WL_TK_ACT[379] WL_TK_ACT[380] 
+ WL_TK_ACT[381] WL_TK_ACT[382] WL_TK_ACT[383] WL_TK_ACT[384] WL_TK_ACT[385] 
+ WL_TK_ACT[386] WL_TK_ACT[387] WL_TK_ACT[388] WL_TK_ACT[389] WL_TK_ACT[390] 
+ WL_TK_ACT[391] WL_TK_ACT[392] WL_TK_ACT[393] WL_TK_ACT[394] WL_TK_ACT[395] 
+ WL_TK_ACT[396] WL_TK_ACT[397] WL_TK_ACT[398] WL_TK_ACT[399] WL_TK_ACT[400] 
+ WL_TK_ACT[401] WL_TK_ACT[402] WL_TK_ACT[403] WL_TK_ACT[404] WL_TK_ACT[405] 
+ WL_TK_ACT[406] WL_TK_ACT[407] WL_TK_ACT[408] WL_TK_ACT[409] WL_TK_ACT[410] 
+ WL_TK_ACT[411] WL_TK_ACT[412] WL_TK_ACT[413] WL_TK_ACT[414] WL_TK_ACT[415] 
+ WL_TK_ACT[416] WL_TK_ACT[417] WL_TK_ACT[418] WL_TK_ACT[419] WL_TK_ACT[420] 
+ WL_TK_ACT[421] WL_TK_ACT[422] WL_TK_ACT[423] WL_TK_ACT[424] WL_TK_ACT[425] 
+ WL_TK_ACT[426] WL_TK_ACT[427] WL_TK_ACT[428] WL_TK_ACT[429] WL_TK_ACT[430] 
+ WL_TK_ACT[431] WL_TK_ACT[432] WL_TK_ACT[433] WL_TK_ACT[434] WL_TK_ACT[435] 
+ WL_TK_ACT[436] WL_TK_ACT[437] WL_TK_ACT[438] WL_TK_ACT[439] WL_TK_ACT[440] 
+ WL_TK_ACT[441] WL_TK_ACT[442] WL_TK_ACT[443] WL_TK_ACT[444] WL_TK_ACT[445] 
+ WL_TK_ACT[446] WL_TK_ACT[447] WL_TK_ACT[448] WL_TK_ACT[449] WL_TK_ACT[450] 
+ WL_TK_ACT[451] WL_TK_ACT[452] WL_TK_ACT[453] WL_TK_ACT[454] WL_TK_ACT[455] 
+ WL_TK_ACT[456] WL_TK_ACT[457] WL_TK_ACT[458] WL_TK_ACT[459] WL_TK_ACT[460] 
+ WL_TK_ACT[461] WL_TK_ACT[462] WL_TK_ACT[463] WL_TK_ACT[464] WL_TK_ACT[465] 
+ WL_TK_ACT[466] WL_TK_ACT[467] WL_TK_ACT[468] WL_TK_ACT[469] WL_TK_ACT[470] 
+ WL_TK_ACT[471] WL_TK_ACT[472] WL_TK_ACT[473] WL_TK_ACT[474] WL_TK_ACT[475] 
+ WL_TK_ACT[476] WL_TK_ACT[477] WL_TK_ACT[478] WL_TK_ACT[479] WL_TK_ACT[480] 
+ WL_TK_ACT[481] WL_TK_ACT[482] WL_TK_ACT[483] WL_TK_ACT[484] WL_TK_ACT[485] 
+ WL_TK_ACT[486] WL_TK_ACT[487] WL_TK_ACT[488] WL_TK_ACT[489] WL_TK_ACT[490] 
+ WL_TK_ACT[491] WL_TK_ACT[492] WL_TK_ACT[493] WL_TK_ACT[494] WL_TK_ACT[495] 
+ WL_TK_ACT[496] WL_TK_ACT[497] WL_TK_ACT[498] WL_TK_ACT[499] WL_TK_ACT[500] 
+ WL_TK_ACT[501] WL_TK_ACT[502] WL_TK_ACT[503] WL_TK_ACT[504] WL_TK_ACT[505] 
+ WL_TK_ACT[506] WL_TK_ACT[507] WL_TK_ACT[508] WL_TK_ACT[509] WL_TK_ACT[510] 
+ WL_TK_ACT[511] TIEH_BT TIEL S1AHSF400W40_TKBL_SIM
XTKWL_LD VDDI TK_R2 TK_R3 VSSI WL_DUM_R2 WL_DUM_R3 WL_TK_R2 WL_TK_R3 
+ S1AHSF400W40_TKWL_LD_SIM
XTKWL_L VDDI TK TK_R2 VSSI WL_DUM_LT WL_DUM_R2 WL_TK WL_TK_R2 S1AHSF400W40_TKWL_SIM
XTKWL_R VDDI TK_R3 NET1095 VSSI WL_DUM_R3 NET939 WL_TK_R3 WL_TK_LD S1AHSF400W40_TKWL_SIM
XIO_RL AWT2_L1 AWT2_R2 BIST2IO_L1 BIST2IO_R2 NET01028 NET01027 CKD_L1 CKD_R2 
+ NET01026 NET01024 NET01023 NET01022 NET01030 NET01029 PD_BUF_1 PD_BUF_R2 
+ NET01025 VDDHD VDDI VSSI WLP_SAEB_L1 WLP_SAEB_R2 S1AHSF400W40_IO_SIM
XIO_LR AWT2_L2 AWT2_L1 BIST2IO_L2 BIST2IO_L1 BWEBM_LR BWEB_LR CKD_L2 CKD_L1 
+ DM_LR D_LR GBLB_LR_12 GBL_LR_12 GWB_LR_12 GW_LR_12 PD_BUF_L2 PD_BUF_1 Q_LR 
+ VDDHD VDDI VSSI WLP_SAEB_L2 WLP_SAEB_L1 S1AHSF400W40_IO_SIM
XIO_LL AWT2_L4 AWT2_L3 BIST2IO_L4 BIST2IO_L3 BWEBM_LL BWEB_LL CKD_L4 CKD_L3 
+ DM_LL D_LL GBLB_LL_12 GBL_LL_12 GWB_LL_12 GW_LL_12 PD_BUF_L4 PD_BUF_L3 Q_LL 
+ VDDHD VDDI VSSI WLP_SAEB_L4 WLP_SAEB_L3 S1AHSF400W40_IO_SIM
XIO_RR AWT2_R3 AWT2_R4 BIST2IO_R3 BIST2IO_R4 NET01006 NET01005 CKD_R3 CKD_R4 
+ NET01004 NET01002 NET01001 NET01000 NET01008 NET01007 PD_BUF_R3 PD_BUF_R4 
+ NET01003 VDDHD VDDI VSSI WLP_SAEB_R3 WLP_SAEB_R4 S1AHSF400W40_IO_SIM
XIO_LD_L AWT2_L3 AWT2_L2 BIST2IO_L3 BIST2IO_L2 CKD_L3 CKD_L2 PD_BUF_L3 
+ PD_BUF_L2 VDDHD VDDI VSSI WLP_SAEB_L3 WLP_SAEB_L2 S1AHSF400W40_IO_LD_SIM
XIO_LD_R AWT2_R2 AWT2_R3 BIST2IO_R2 BIST2IO_R3 CKD_R2 CKD_R3 PD_BUF_R2 
+ PD_BUF_R3 VDDHD VDDI VSSI WLP_SAEB_R2 WLP_SAEB_R3 S1AHSF400W40_IO_LD_SIM
XCNT AWT AWT2_L1 BIST BIST2IO_L1 WL_TK CEB CEBM CKD_L1 CLK VDDHD VDDI 
+ DEC_X0_1[0] DEC_X0_1[1] DEC_X0_1[2] DEC_X0_1[3] DEC_X0_1[4] DEC_X0_1[5] 
+ DEC_X0_1[6] DEC_X0_1[7] DEC_X1_1[0] DEC_X1_1[1] DEC_X1_1[2] DEC_X1_1[3] 
+ DEC_X1_1[4] DEC_X1_1[5] DEC_X1_1[6] DEC_X1_1[7] DEC_X2_1[0] DEC_X2_1[1] 
+ DEC_X2_1[2] DEC_X2_1[3] DEC_X3_1[0] DEC_X3_1[1] DEC_X3_1[2] DEC_X3_1[3] 
+ DEC_X3_1[4] DEC_X3_1[5] DEC_X3_1[6] DEC_X3_1[7] DEC_Y_1[0] DEC_Y_1[1] 
+ DEC_Y_1[2] DEC_Y_1[3] DEC_Y_1[4] DEC_Y_1[5] DEC_Y_1[6] DEC_Y_1[7] FAD1[0] 
+ FAD1[1] FAD1[2] FAD1[3] FAD1[4] FAD1[5] FAD1[6] FAD1[7] FAD1[8] FAD1[9] 
+ FAD1[10] FAD2[0] FAD2[1] FAD2[2] FAD2[3] FAD2[4] FAD2[5] FAD2[6] FAD2[7] 
+ FAD2[8] FAD2[9] FAD2[10] NET1083[0] NET1083[1] PD PD_BUF_1 PD_CVDDBUF_1 
+ PTSEL REDEN_BT REDEN1 REDEN2 REDENB_BT RSTB RTSEL[0] RTSEL[1] RW_RE_1 SCLK 
+ SDIN SDOUT TK TM TRKBL VDDHD VDDI VHI_LT VLO_LT VSSI WEB WEBM WLP_SAE_1 
+ WLP_SAEB_L1 WLP_SAE_TK_1 WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] 
+ X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] 
+ XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL_1[0] YM[0] YM[1] YM[2] YM[3] 
+ S1AHSF400W40_CNT_SIM
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    SIM_ALL
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_SIM_ALL
*.PININFO
XI7 NET075 NET074 NET073 NET068 NET067 NET060 NET071 NET070 NET069 NET059 
+ NET058 NET057 NET056 NET066 NET080 NET079 NET076 NET077[0] NET077[1] NET063 
+ NET053 NET052 NET062 NET061 NET088[0] NET088[1] NET088[2] NET088[3] 
+ NET088[4] NET088[5] NET088[6] NET088[7] NET088[8] NET088[9] NET088[10] 
+ NET088[11] NET088[12] NET088[13] NET088[14] NET088[15] NET088[16] NET088[17] 
+ NET088[18] NET088[19] NET088[20] NET088[21] NET088[22] NET088[23] NET088[24] 
+ NET088[25] NET088[26] NET088[27] NET088[28] NET088[29] NET088[30] NET088[31] 
+ NET088[32] NET088[33] NET088[34] NET088[35] NET088[36] NET088[37] NET088[38] 
+ NET088[39] NET088[40] NET088[41] NET088[42] NET088[43] NET088[44] NET088[45] 
+ NET088[46] NET088[47] NET088[48] NET088[49] NET088[50] NET088[51] NET088[52] 
+ NET088[53] NET088[54] NET088[55] NET088[56] NET088[57] NET088[58] NET088[59] 
+ NET088[60] NET088[61] NET088[62] NET088[63] NET088[64] NET088[65] NET088[66] 
+ NET088[67] NET088[68] NET088[69] NET088[70] NET088[71] NET088[72] NET088[73] 
+ NET088[74] NET088[75] NET088[76] NET088[77] NET088[78] NET088[79] NET088[80] 
+ NET088[81] NET088[82] NET088[83] NET088[84] NET088[85] NET088[86] NET088[87] 
+ NET088[88] NET088[89] NET088[90] NET088[91] NET088[92] NET088[93] NET088[94] 
+ NET088[95] NET088[96] NET088[97] NET088[98] NET088[99] NET088[100] 
+ NET088[101] NET088[102] NET088[103] NET088[104] NET088[105] NET088[106] 
+ NET088[107] NET088[108] NET088[109] NET088[110] NET088[111] NET088[112] 
+ NET088[113] NET088[114] NET088[115] NET088[116] NET088[117] NET088[118] 
+ NET088[119] NET088[120] NET088[121] NET088[122] NET088[123] NET088[124] 
+ NET088[125] NET088[126] NET088[127] NET088[128] NET088[129] NET088[130] 
+ NET088[131] NET088[132] NET088[133] NET088[134] NET088[135] NET088[136] 
+ NET088[137] NET088[138] NET088[139] NET088[140] NET088[141] NET088[142] 
+ NET088[143] NET088[144] NET088[145] NET088[146] NET088[147] NET088[148] 
+ NET088[149] NET088[150] NET088[151] NET088[152] NET088[153] NET088[154] 
+ NET088[155] NET088[156] NET088[157] NET088[158] NET088[159] NET088[160] 
+ NET088[161] NET088[162] NET088[163] NET088[164] NET088[165] NET088[166] 
+ NET088[167] NET088[168] NET088[169] NET088[170] NET088[171] NET088[172] 
+ NET088[173] NET088[174] NET088[175] NET088[176] NET088[177] NET088[178] 
+ NET088[179] NET088[180] NET088[181] NET088[182] NET088[183] NET088[184] 
+ NET088[185] NET088[186] NET088[187] NET088[188] NET088[189] NET088[190] 
+ NET088[191] NET088[192] NET088[193] NET088[194] NET088[195] NET088[196] 
+ NET088[197] NET088[198] NET088[199] NET088[200] NET088[201] NET088[202] 
+ NET088[203] NET088[204] NET088[205] NET088[206] NET088[207] NET088[208] 
+ NET088[209] NET088[210] NET088[211] NET088[212] NET088[213] NET088[214] 
+ NET088[215] NET088[216] NET088[217] NET088[218] NET088[219] NET088[220] 
+ NET088[221] NET088[222] NET088[223] NET088[224] NET088[225] NET088[226] 
+ NET088[227] NET088[228] NET088[229] NET088[230] NET088[231] NET088[232] 
+ NET088[233] NET088[234] NET088[235] NET088[236] NET088[237] NET088[238] 
+ NET088[239] NET088[240] NET088[241] NET088[242] NET088[243] NET088[244] 
+ NET088[245] NET088[246] NET088[247] NET088[248] NET088[249] NET088[250] 
+ NET088[251] NET088[252] NET088[253] NET088[254] NET088[255] NET088[256] 
+ NET088[257] NET088[258] NET088[259] NET088[260] NET088[261] NET088[262] 
+ NET088[263] NET088[264] NET088[265] NET088[266] NET088[267] NET088[268] 
+ NET088[269] NET088[270] NET088[271] NET088[272] NET088[273] NET088[274] 
+ NET088[275] NET088[276] NET088[277] NET088[278] NET088[279] NET088[280] 
+ NET088[281] NET088[282] NET088[283] NET088[284] NET088[285] NET088[286] 
+ NET088[287] NET088[288] NET088[289] NET088[290] NET088[291] NET088[292] 
+ NET088[293] NET088[294] NET088[295] NET088[296] NET088[297] NET088[298] 
+ NET088[299] NET088[300] NET088[301] NET088[302] NET088[303] NET088[304] 
+ NET088[305] NET088[306] NET088[307] NET088[308] NET088[309] NET088[310] 
+ NET088[311] NET088[312] NET088[313] NET088[314] NET088[315] NET088[316] 
+ NET088[317] NET088[318] NET088[319] NET088[320] NET088[321] NET088[322] 
+ NET088[323] NET088[324] NET088[325] NET088[326] NET088[327] NET088[328] 
+ NET088[329] NET088[330] NET088[331] NET088[332] NET088[333] NET088[334] 
+ NET088[335] NET088[336] NET088[337] NET088[338] NET088[339] NET088[340] 
+ NET088[341] NET088[342] NET088[343] NET088[344] NET088[345] NET088[346] 
+ NET088[347] NET088[348] NET088[349] NET088[350] NET088[351] NET088[352] 
+ NET088[353] NET088[354] NET088[355] NET088[356] NET088[357] NET088[358] 
+ NET088[359] NET088[360] NET088[361] NET088[362] NET088[363] NET088[364] 
+ NET088[365] NET088[366] NET088[367] NET088[368] NET088[369] NET088[370] 
+ NET088[371] NET088[372] NET088[373] NET088[374] NET088[375] NET088[376] 
+ NET088[377] NET088[378] NET088[379] NET088[380] NET088[381] NET088[382] 
+ NET088[383] NET088[384] NET088[385] NET088[386] NET088[387] NET088[388] 
+ NET088[389] NET088[390] NET088[391] NET088[392] NET088[393] NET088[394] 
+ NET088[395] NET088[396] NET088[397] NET088[398] NET088[399] NET088[400] 
+ NET088[401] NET088[402] NET088[403] NET088[404] NET088[405] NET088[406] 
+ NET088[407] NET088[408] NET088[409] NET088[410] NET088[411] NET088[412] 
+ NET088[413] NET088[414] NET088[415] NET088[416] NET088[417] NET088[418] 
+ NET088[419] NET088[420] NET088[421] NET088[422] NET088[423] NET088[424] 
+ NET088[425] NET088[426] NET088[427] NET088[428] NET088[429] NET088[430] 
+ NET088[431] NET088[432] NET088[433] NET088[434] NET088[435] NET088[436] 
+ NET088[437] NET088[438] NET088[439] NET088[440] NET088[441] NET088[442] 
+ NET088[443] NET088[444] NET088[445] NET088[446] NET088[447] NET088[448] 
+ NET088[449] NET088[450] NET088[451] NET088[452] NET088[453] NET088[454] 
+ NET088[455] NET088[456] NET088[457] NET088[458] NET088[459] NET088[460] 
+ NET088[461] NET088[462] NET088[463] NET088[464] NET088[465] NET088[466] 
+ NET088[467] NET088[468] NET088[469] NET088[470] NET088[471] NET088[472] 
+ NET088[473] NET088[474] NET088[475] NET088[476] NET088[477] NET088[478] 
+ NET088[479] NET088[480] NET088[481] NET088[482] NET088[483] NET088[484] 
+ NET088[485] NET088[486] NET088[487] NET088[488] NET088[489] NET088[490] 
+ NET088[491] NET088[492] NET088[493] NET088[494] NET088[495] NET088[496] 
+ NET088[497] NET088[498] NET088[499] NET088[500] NET088[501] NET088[502] 
+ NET088[503] NET088[504] NET088[505] NET088[506] NET088[507] NET088[508] 
+ NET088[509] NET088[510] NET088[511] NET078 NET072[0] NET072[1] NET072[2] 
+ NET065[0] NET065[1] NET065[2] NET065[3] NET065[4] NET065[5] NET065[6] 
+ NET065[7] NET065[8] NET064[0] NET064[1] NET064[2] NET064[3] NET064[4] 
+ NET064[5] NET064[6] NET064[7] NET064[8] NET055[0] NET055[1] NET055[2] 
+ NET055[3] NET054[0] NET054[1] NET054[2] NET054[3] S1AHSF400W40_SIM_SB1S
XI6 NET0138 NET0137 NET0135 NET0131 NET0130 NET0117 NET0134 NET0133 NET0132 
+ NET0116 NET0115 NET0114 NET0113 NET0146[0] NET0146[1] NET0146[2] NET0146[3] 
+ NET0146[4] NET0146[5] NET0146[6] NET0146[7] NET0146[8] NET0146[9] 
+ NET0146[10] NET0145[0] NET0145[1] NET0145[2] NET0145[3] NET0145[4] 
+ NET0145[5] NET0145[6] NET0145[7] NET0145[8] NET0145[9] NET0145[10] NET0128 
+ NET0127 NET0142 NET0140 NET0126 NET0125 NET0124 NET0144[0] NET0144[1] 
+ NET0122 NET0121 NET0139 NET0120 NET040 NET039 NET0119 NET0118 NET045[0] 
+ NET045[1] NET045[2] NET045[3] NET045[4] NET045[5] NET045[6] NET045[7] 
+ NET045[8] NET045[9] NET045[10] NET045[11] NET045[12] NET045[13] NET045[14] 
+ NET045[15] NET045[16] NET045[17] NET045[18] NET045[19] NET045[20] NET045[21] 
+ NET045[22] NET045[23] NET045[24] NET045[25] NET045[26] NET045[27] NET045[28] 
+ NET045[29] NET045[30] NET045[31] NET045[32] NET045[33] NET045[34] NET045[35] 
+ NET045[36] NET045[37] NET045[38] NET045[39] NET045[40] NET045[41] NET045[42] 
+ NET045[43] NET045[44] NET045[45] NET045[46] NET045[47] NET045[48] NET045[49] 
+ NET045[50] NET045[51] NET045[52] NET045[53] NET045[54] NET045[55] NET045[56] 
+ NET045[57] NET045[58] NET045[59] NET045[60] NET045[61] NET045[62] NET045[63] 
+ NET045[64] NET045[65] NET045[66] NET045[67] NET045[68] NET045[69] NET045[70] 
+ NET045[71] NET045[72] NET045[73] NET045[74] NET045[75] NET045[76] NET045[77] 
+ NET045[78] NET045[79] NET045[80] NET045[81] NET045[82] NET045[83] NET045[84] 
+ NET045[85] NET045[86] NET045[87] NET045[88] NET045[89] NET045[90] NET045[91] 
+ NET045[92] NET045[93] NET045[94] NET045[95] NET045[96] NET045[97] NET045[98] 
+ NET045[99] NET045[100] NET045[101] NET045[102] NET045[103] NET045[104] 
+ NET045[105] NET045[106] NET045[107] NET045[108] NET045[109] NET045[110] 
+ NET045[111] NET045[112] NET045[113] NET045[114] NET045[115] NET045[116] 
+ NET045[117] NET045[118] NET045[119] NET045[120] NET045[121] NET045[122] 
+ NET045[123] NET045[124] NET045[125] NET045[126] NET045[127] NET045[128] 
+ NET045[129] NET045[130] NET045[131] NET045[132] NET045[133] NET045[134] 
+ NET045[135] NET045[136] NET045[137] NET045[138] NET045[139] NET045[140] 
+ NET045[141] NET045[142] NET045[143] NET045[144] NET045[145] NET045[146] 
+ NET045[147] NET045[148] NET045[149] NET045[150] NET045[151] NET045[152] 
+ NET045[153] NET045[154] NET045[155] NET045[156] NET045[157] NET045[158] 
+ NET045[159] NET045[160] NET045[161] NET045[162] NET045[163] NET045[164] 
+ NET045[165] NET045[166] NET045[167] NET045[168] NET045[169] NET045[170] 
+ NET045[171] NET045[172] NET045[173] NET045[174] NET045[175] NET045[176] 
+ NET045[177] NET045[178] NET045[179] NET045[180] NET045[181] NET045[182] 
+ NET045[183] NET045[184] NET045[185] NET045[186] NET045[187] NET045[188] 
+ NET045[189] NET045[190] NET045[191] NET045[192] NET045[193] NET045[194] 
+ NET045[195] NET045[196] NET045[197] NET045[198] NET045[199] NET045[200] 
+ NET045[201] NET045[202] NET045[203] NET045[204] NET045[205] NET045[206] 
+ NET045[207] NET045[208] NET045[209] NET045[210] NET045[211] NET045[212] 
+ NET045[213] NET045[214] NET045[215] NET045[216] NET045[217] NET045[218] 
+ NET045[219] NET045[220] NET045[221] NET045[222] NET045[223] NET045[224] 
+ NET045[225] NET045[226] NET045[227] NET045[228] NET045[229] NET045[230] 
+ NET045[231] NET045[232] NET045[233] NET045[234] NET045[235] NET045[236] 
+ NET045[237] NET045[238] NET045[239] NET045[240] NET045[241] NET045[242] 
+ NET045[243] NET045[244] NET045[245] NET045[246] NET045[247] NET045[248] 
+ NET045[249] NET045[250] NET045[251] NET045[252] NET045[253] NET045[254] 
+ NET045[255] NET045[256] NET045[257] NET045[258] NET045[259] NET045[260] 
+ NET045[261] NET045[262] NET045[263] NET045[264] NET045[265] NET045[266] 
+ NET045[267] NET045[268] NET045[269] NET045[270] NET045[271] NET045[272] 
+ NET045[273] NET045[274] NET045[275] NET045[276] NET045[277] NET045[278] 
+ NET045[279] NET045[280] NET045[281] NET045[282] NET045[283] NET045[284] 
+ NET045[285] NET045[286] NET045[287] NET045[288] NET045[289] NET045[290] 
+ NET045[291] NET045[292] NET045[293] NET045[294] NET045[295] NET045[296] 
+ NET045[297] NET045[298] NET045[299] NET045[300] NET045[301] NET045[302] 
+ NET045[303] NET045[304] NET045[305] NET045[306] NET045[307] NET045[308] 
+ NET045[309] NET045[310] NET045[311] NET045[312] NET045[313] NET045[314] 
+ NET045[315] NET045[316] NET045[317] NET045[318] NET045[319] NET045[320] 
+ NET045[321] NET045[322] NET045[323] NET045[324] NET045[325] NET045[326] 
+ NET045[327] NET045[328] NET045[329] NET045[330] NET045[331] NET045[332] 
+ NET045[333] NET045[334] NET045[335] NET045[336] NET045[337] NET045[338] 
+ NET045[339] NET045[340] NET045[341] NET045[342] NET045[343] NET045[344] 
+ NET045[345] NET045[346] NET045[347] NET045[348] NET045[349] NET045[350] 
+ NET045[351] NET045[352] NET045[353] NET045[354] NET045[355] NET045[356] 
+ NET045[357] NET045[358] NET045[359] NET045[360] NET045[361] NET045[362] 
+ NET045[363] NET045[364] NET045[365] NET045[366] NET045[367] NET045[368] 
+ NET045[369] NET045[370] NET045[371] NET045[372] NET045[373] NET045[374] 
+ NET045[375] NET045[376] NET045[377] NET045[378] NET045[379] NET045[380] 
+ NET045[381] NET045[382] NET045[383] NET045[384] NET045[385] NET045[386] 
+ NET045[387] NET045[388] NET045[389] NET045[390] NET045[391] NET045[392] 
+ NET045[393] NET045[394] NET045[395] NET045[396] NET045[397] NET045[398] 
+ NET045[399] NET045[400] NET045[401] NET045[402] NET045[403] NET045[404] 
+ NET045[405] NET045[406] NET045[407] NET045[408] NET045[409] NET045[410] 
+ NET045[411] NET045[412] NET045[413] NET045[414] NET045[415] NET045[416] 
+ NET045[417] NET045[418] NET045[419] NET045[420] NET045[421] NET045[422] 
+ NET045[423] NET045[424] NET045[425] NET045[426] NET045[427] NET045[428] 
+ NET045[429] NET045[430] NET045[431] NET045[432] NET045[433] NET045[434] 
+ NET045[435] NET045[436] NET045[437] NET045[438] NET045[439] NET045[440] 
+ NET045[441] NET045[442] NET045[443] NET045[444] NET045[445] NET045[446] 
+ NET045[447] NET045[448] NET045[449] NET045[450] NET045[451] NET045[452] 
+ NET045[453] NET045[454] NET045[455] NET045[456] NET045[457] NET045[458] 
+ NET045[459] NET045[460] NET045[461] NET045[462] NET045[463] NET045[464] 
+ NET045[465] NET045[466] NET045[467] NET045[468] NET045[469] NET045[470] 
+ NET045[471] NET045[472] NET045[473] NET045[474] NET045[475] NET045[476] 
+ NET045[477] NET045[478] NET045[479] NET045[480] NET045[481] NET045[482] 
+ NET045[483] NET045[484] NET045[485] NET045[486] NET045[487] NET045[488] 
+ NET045[489] NET045[490] NET045[491] NET045[492] NET045[493] NET045[494] 
+ NET045[495] NET045[496] NET045[497] NET045[498] NET045[499] NET045[500] 
+ NET045[501] NET045[502] NET045[503] NET045[504] NET045[505] NET045[506] 
+ NET045[507] NET045[508] NET045[509] NET045[510] NET045[511] NET0143 
+ NET0136[0] NET0136[1] NET0136[2] NET0129[0] NET0129[1] NET0129[2] NET0129[3] 
+ NET0129[4] NET0129[5] NET0129[6] NET0129[7] NET0129[8] NET0129[9] 
+ NET0129[10] NET0123[0] NET0123[1] NET0123[2] NET0123[3] NET0123[4] 
+ NET0123[5] NET0123[6] NET0123[7] NET0123[8] NET0123[9] NET0123[10] 
+ NET0112[0] NET0112[1] NET0112[2] NET0112[3] NET0111[0] NET0111[1] NET0111[2] 
+ NET0111[3] S1AHSF400W40_SIM_HB
XI5 NET030 NET029 NET027 NET023 NET022 NET09 NET026 NET025 NET024 NET08 NET07 
+ NET06 NET05 NET038[0] NET038[1] NET038[2] NET038[3] NET038[4] NET038[5] 
+ NET038[6] NET038[7] NET038[8] NET038[9] NET038[10] NET037[0] NET037[1] 
+ NET037[2] NET037[3] NET037[4] NET037[5] NET037[6] NET037[7] NET037[8] 
+ NET037[9] NET037[10] NET020 NET019 NET034 NET0107 NET018 NET017 NET016 
+ NET036[0] NET036[1] NET014 NET013 NET0109 NET012 NET0110 NET0108 NET011 
+ NET010 NET0156[0] NET0156[1] NET0156[2] NET0156[3] NET0156[4] NET0156[5] 
+ NET0156[6] NET0156[7] NET0156[8] NET0156[9] NET0156[10] NET0156[11] 
+ NET0156[12] NET0156[13] NET0156[14] NET0156[15] NET0156[16] NET0156[17] 
+ NET0156[18] NET0156[19] NET0156[20] NET0156[21] NET0156[22] NET0156[23] 
+ NET0156[24] NET0156[25] NET0156[26] NET0156[27] NET0156[28] NET0156[29] 
+ NET0156[30] NET0156[31] NET0156[32] NET0156[33] NET0156[34] NET0156[35] 
+ NET0156[36] NET0156[37] NET0156[38] NET0156[39] NET0156[40] NET0156[41] 
+ NET0156[42] NET0156[43] NET0156[44] NET0156[45] NET0156[46] NET0156[47] 
+ NET0156[48] NET0156[49] NET0156[50] NET0156[51] NET0156[52] NET0156[53] 
+ NET0156[54] NET0156[55] NET0156[56] NET0156[57] NET0156[58] NET0156[59] 
+ NET0156[60] NET0156[61] NET0156[62] NET0156[63] NET0156[64] NET0156[65] 
+ NET0156[66] NET0156[67] NET0156[68] NET0156[69] NET0156[70] NET0156[71] 
+ NET0156[72] NET0156[73] NET0156[74] NET0156[75] NET0156[76] NET0156[77] 
+ NET0156[78] NET0156[79] NET0156[80] NET0156[81] NET0156[82] NET0156[83] 
+ NET0156[84] NET0156[85] NET0156[86] NET0156[87] NET0156[88] NET0156[89] 
+ NET0156[90] NET0156[91] NET0156[92] NET0156[93] NET0156[94] NET0156[95] 
+ NET0156[96] NET0156[97] NET0156[98] NET0156[99] NET0156[100] NET0156[101] 
+ NET0156[102] NET0156[103] NET0156[104] NET0156[105] NET0156[106] 
+ NET0156[107] NET0156[108] NET0156[109] NET0156[110] NET0156[111] 
+ NET0156[112] NET0156[113] NET0156[114] NET0156[115] NET0156[116] 
+ NET0156[117] NET0156[118] NET0156[119] NET0156[120] NET0156[121] 
+ NET0156[122] NET0156[123] NET0156[124] NET0156[125] NET0156[126] 
+ NET0156[127] NET0156[128] NET0156[129] NET0156[130] NET0156[131] 
+ NET0156[132] NET0156[133] NET0156[134] NET0156[135] NET0156[136] 
+ NET0156[137] NET0156[138] NET0156[139] NET0156[140] NET0156[141] 
+ NET0156[142] NET0156[143] NET0156[144] NET0156[145] NET0156[146] 
+ NET0156[147] NET0156[148] NET0156[149] NET0156[150] NET0156[151] 
+ NET0156[152] NET0156[153] NET0156[154] NET0156[155] NET0156[156] 
+ NET0156[157] NET0156[158] NET0156[159] NET0156[160] NET0156[161] 
+ NET0156[162] NET0156[163] NET0156[164] NET0156[165] NET0156[166] 
+ NET0156[167] NET0156[168] NET0156[169] NET0156[170] NET0156[171] 
+ NET0156[172] NET0156[173] NET0156[174] NET0156[175] NET0156[176] 
+ NET0156[177] NET0156[178] NET0156[179] NET0156[180] NET0156[181] 
+ NET0156[182] NET0156[183] NET0156[184] NET0156[185] NET0156[186] 
+ NET0156[187] NET0156[188] NET0156[189] NET0156[190] NET0156[191] 
+ NET0156[192] NET0156[193] NET0156[194] NET0156[195] NET0156[196] 
+ NET0156[197] NET0156[198] NET0156[199] NET0156[200] NET0156[201] 
+ NET0156[202] NET0156[203] NET0156[204] NET0156[205] NET0156[206] 
+ NET0156[207] NET0156[208] NET0156[209] NET0156[210] NET0156[211] 
+ NET0156[212] NET0156[213] NET0156[214] NET0156[215] NET0156[216] 
+ NET0156[217] NET0156[218] NET0156[219] NET0156[220] NET0156[221] 
+ NET0156[222] NET0156[223] NET0156[224] NET0156[225] NET0156[226] 
+ NET0156[227] NET0156[228] NET0156[229] NET0156[230] NET0156[231] 
+ NET0156[232] NET0156[233] NET0156[234] NET0156[235] NET0156[236] 
+ NET0156[237] NET0156[238] NET0156[239] NET0156[240] NET0156[241] 
+ NET0156[242] NET0156[243] NET0156[244] NET0156[245] NET0156[246] 
+ NET0156[247] NET0156[248] NET0156[249] NET0156[250] NET0156[251] 
+ NET0156[252] NET0156[253] NET0156[254] NET0156[255] NET0156[256] 
+ NET0156[257] NET0156[258] NET0156[259] NET0156[260] NET0156[261] 
+ NET0156[262] NET0156[263] NET0156[264] NET0156[265] NET0156[266] 
+ NET0156[267] NET0156[268] NET0156[269] NET0156[270] NET0156[271] 
+ NET0156[272] NET0156[273] NET0156[274] NET0156[275] NET0156[276] 
+ NET0156[277] NET0156[278] NET0156[279] NET0156[280] NET0156[281] 
+ NET0156[282] NET0156[283] NET0156[284] NET0156[285] NET0156[286] 
+ NET0156[287] NET0156[288] NET0156[289] NET0156[290] NET0156[291] 
+ NET0156[292] NET0156[293] NET0156[294] NET0156[295] NET0156[296] 
+ NET0156[297] NET0156[298] NET0156[299] NET0156[300] NET0156[301] 
+ NET0156[302] NET0156[303] NET0156[304] NET0156[305] NET0156[306] 
+ NET0156[307] NET0156[308] NET0156[309] NET0156[310] NET0156[311] 
+ NET0156[312] NET0156[313] NET0156[314] NET0156[315] NET0156[316] 
+ NET0156[317] NET0156[318] NET0156[319] NET0156[320] NET0156[321] 
+ NET0156[322] NET0156[323] NET0156[324] NET0156[325] NET0156[326] 
+ NET0156[327] NET0156[328] NET0156[329] NET0156[330] NET0156[331] 
+ NET0156[332] NET0156[333] NET0156[334] NET0156[335] NET0156[336] 
+ NET0156[337] NET0156[338] NET0156[339] NET0156[340] NET0156[341] 
+ NET0156[342] NET0156[343] NET0156[344] NET0156[345] NET0156[346] 
+ NET0156[347] NET0156[348] NET0156[349] NET0156[350] NET0156[351] 
+ NET0156[352] NET0156[353] NET0156[354] NET0156[355] NET0156[356] 
+ NET0156[357] NET0156[358] NET0156[359] NET0156[360] NET0156[361] 
+ NET0156[362] NET0156[363] NET0156[364] NET0156[365] NET0156[366] 
+ NET0156[367] NET0156[368] NET0156[369] NET0156[370] NET0156[371] 
+ NET0156[372] NET0156[373] NET0156[374] NET0156[375] NET0156[376] 
+ NET0156[377] NET0156[378] NET0156[379] NET0156[380] NET0156[381] 
+ NET0156[382] NET0156[383] NET0156[384] NET0156[385] NET0156[386] 
+ NET0156[387] NET0156[388] NET0156[389] NET0156[390] NET0156[391] 
+ NET0156[392] NET0156[393] NET0156[394] NET0156[395] NET0156[396] 
+ NET0156[397] NET0156[398] NET0156[399] NET0156[400] NET0156[401] 
+ NET0156[402] NET0156[403] NET0156[404] NET0156[405] NET0156[406] 
+ NET0156[407] NET0156[408] NET0156[409] NET0156[410] NET0156[411] 
+ NET0156[412] NET0156[413] NET0156[414] NET0156[415] NET0156[416] 
+ NET0156[417] NET0156[418] NET0156[419] NET0156[420] NET0156[421] 
+ NET0156[422] NET0156[423] NET0156[424] NET0156[425] NET0156[426] 
+ NET0156[427] NET0156[428] NET0156[429] NET0156[430] NET0156[431] 
+ NET0156[432] NET0156[433] NET0156[434] NET0156[435] NET0156[436] 
+ NET0156[437] NET0156[438] NET0156[439] NET0156[440] NET0156[441] 
+ NET0156[442] NET0156[443] NET0156[444] NET0156[445] NET0156[446] 
+ NET0156[447] NET0156[448] NET0156[449] NET0156[450] NET0156[451] 
+ NET0156[452] NET0156[453] NET0156[454] NET0156[455] NET0156[456] 
+ NET0156[457] NET0156[458] NET0156[459] NET0156[460] NET0156[461] 
+ NET0156[462] NET0156[463] NET0156[464] NET0156[465] NET0156[466] 
+ NET0156[467] NET0156[468] NET0156[469] NET0156[470] NET0156[471] 
+ NET0156[472] NET0156[473] NET0156[474] NET0156[475] NET0156[476] 
+ NET0156[477] NET0156[478] NET0156[479] NET0156[480] NET0156[481] 
+ NET0156[482] NET0156[483] NET0156[484] NET0156[485] NET0156[486] 
+ NET0156[487] NET0156[488] NET0156[489] NET0156[490] NET0156[491] 
+ NET0156[492] NET0156[493] NET0156[494] NET0156[495] NET0156[496] 
+ NET0156[497] NET0156[498] NET0156[499] NET0156[500] NET0156[501] 
+ NET0156[502] NET0156[503] NET0156[504] NET0156[505] NET0156[506] 
+ NET0156[507] NET0156[508] NET0156[509] NET0156[510] NET0156[511] NET035 
+ NET028[0] NET028[1] NET028[2] NET021[0] NET021[1] NET021[2] NET021[3] 
+ NET021[4] NET021[5] NET021[6] NET021[7] NET021[8] NET021[9] NET021[10] 
+ NET015[0] NET015[1] NET015[2] NET015[3] NET015[4] NET015[5] NET015[6] 
+ NET015[7] NET015[8] NET015[9] NET015[10] NET04[0] NET04[1] NET04[2] NET04[3] 
+ NET03[0] NET03[1] NET03[2] NET03[3] S1AHSF400W40_SIM_1B
XI4 NET24 NET23 NET22 NET17 NET16 NET9 NET20 NET19 NET18 NET8 NET7 NET6 NET5 
+ NET15 NET28 NET27 NET25 NET26[0] NET26[1] NET12 NET2 NET1 NET11 NET10 
+ NET0194[0] NET0194[1] NET0194[2] NET0194[3] NET0194[4] NET0194[5] NET0194[6] 
+ NET0194[7] NET0194[8] NET0194[9] NET0194[10] NET0194[11] NET0194[12] 
+ NET0194[13] NET0194[14] NET0194[15] NET0194[16] NET0194[17] NET0194[18] 
+ NET0194[19] NET0194[20] NET0194[21] NET0194[22] NET0194[23] NET0194[24] 
+ NET0194[25] NET0194[26] NET0194[27] NET0194[28] NET0194[29] NET0194[30] 
+ NET0194[31] NET0194[32] NET0194[33] NET0194[34] NET0194[35] NET0194[36] 
+ NET0194[37] NET0194[38] NET0194[39] NET0194[40] NET0194[41] NET0194[42] 
+ NET0194[43] NET0194[44] NET0194[45] NET0194[46] NET0194[47] NET0194[48] 
+ NET0194[49] NET0194[50] NET0194[51] NET0194[52] NET0194[53] NET0194[54] 
+ NET0194[55] NET0194[56] NET0194[57] NET0194[58] NET0194[59] NET0194[60] 
+ NET0194[61] NET0194[62] NET0194[63] NET0194[64] NET0194[65] NET0194[66] 
+ NET0194[67] NET0194[68] NET0194[69] NET0194[70] NET0194[71] NET0194[72] 
+ NET0194[73] NET0194[74] NET0194[75] NET0194[76] NET0194[77] NET0194[78] 
+ NET0194[79] NET0194[80] NET0194[81] NET0194[82] NET0194[83] NET0194[84] 
+ NET0194[85] NET0194[86] NET0194[87] NET0194[88] NET0194[89] NET0194[90] 
+ NET0194[91] NET0194[92] NET0194[93] NET0194[94] NET0194[95] NET0194[96] 
+ NET0194[97] NET0194[98] NET0194[99] NET0194[100] NET0194[101] NET0194[102] 
+ NET0194[103] NET0194[104] NET0194[105] NET0194[106] NET0194[107] 
+ NET0194[108] NET0194[109] NET0194[110] NET0194[111] NET0194[112] 
+ NET0194[113] NET0194[114] NET0194[115] NET0194[116] NET0194[117] 
+ NET0194[118] NET0194[119] NET0194[120] NET0194[121] NET0194[122] 
+ NET0194[123] NET0194[124] NET0194[125] NET0194[126] NET0194[127] 
+ NET0194[128] NET0194[129] NET0194[130] NET0194[131] NET0194[132] 
+ NET0194[133] NET0194[134] NET0194[135] NET0194[136] NET0194[137] 
+ NET0194[138] NET0194[139] NET0194[140] NET0194[141] NET0194[142] 
+ NET0194[143] NET0194[144] NET0194[145] NET0194[146] NET0194[147] 
+ NET0194[148] NET0194[149] NET0194[150] NET0194[151] NET0194[152] 
+ NET0194[153] NET0194[154] NET0194[155] NET0194[156] NET0194[157] 
+ NET0194[158] NET0194[159] NET0194[160] NET0194[161] NET0194[162] 
+ NET0194[163] NET0194[164] NET0194[165] NET0194[166] NET0194[167] 
+ NET0194[168] NET0194[169] NET0194[170] NET0194[171] NET0194[172] 
+ NET0194[173] NET0194[174] NET0194[175] NET0194[176] NET0194[177] 
+ NET0194[178] NET0194[179] NET0194[180] NET0194[181] NET0194[182] 
+ NET0194[183] NET0194[184] NET0194[185] NET0194[186] NET0194[187] 
+ NET0194[188] NET0194[189] NET0194[190] NET0194[191] NET0194[192] 
+ NET0194[193] NET0194[194] NET0194[195] NET0194[196] NET0194[197] 
+ NET0194[198] NET0194[199] NET0194[200] NET0194[201] NET0194[202] 
+ NET0194[203] NET0194[204] NET0194[205] NET0194[206] NET0194[207] 
+ NET0194[208] NET0194[209] NET0194[210] NET0194[211] NET0194[212] 
+ NET0194[213] NET0194[214] NET0194[215] NET0194[216] NET0194[217] 
+ NET0194[218] NET0194[219] NET0194[220] NET0194[221] NET0194[222] 
+ NET0194[223] NET0194[224] NET0194[225] NET0194[226] NET0194[227] 
+ NET0194[228] NET0194[229] NET0194[230] NET0194[231] NET0194[232] 
+ NET0194[233] NET0194[234] NET0194[235] NET0194[236] NET0194[237] 
+ NET0194[238] NET0194[239] NET0194[240] NET0194[241] NET0194[242] 
+ NET0194[243] NET0194[244] NET0194[245] NET0194[246] NET0194[247] 
+ NET0194[248] NET0194[249] NET0194[250] NET0194[251] NET0194[252] 
+ NET0194[253] NET0194[254] NET0194[255] NET0194[256] NET0194[257] 
+ NET0194[258] NET0194[259] NET0194[260] NET0194[261] NET0194[262] 
+ NET0194[263] NET0194[264] NET0194[265] NET0194[266] NET0194[267] 
+ NET0194[268] NET0194[269] NET0194[270] NET0194[271] NET0194[272] 
+ NET0194[273] NET0194[274] NET0194[275] NET0194[276] NET0194[277] 
+ NET0194[278] NET0194[279] NET0194[280] NET0194[281] NET0194[282] 
+ NET0194[283] NET0194[284] NET0194[285] NET0194[286] NET0194[287] 
+ NET0194[288] NET0194[289] NET0194[290] NET0194[291] NET0194[292] 
+ NET0194[293] NET0194[294] NET0194[295] NET0194[296] NET0194[297] 
+ NET0194[298] NET0194[299] NET0194[300] NET0194[301] NET0194[302] 
+ NET0194[303] NET0194[304] NET0194[305] NET0194[306] NET0194[307] 
+ NET0194[308] NET0194[309] NET0194[310] NET0194[311] NET0194[312] 
+ NET0194[313] NET0194[314] NET0194[315] NET0194[316] NET0194[317] 
+ NET0194[318] NET0194[319] NET0194[320] NET0194[321] NET0194[322] 
+ NET0194[323] NET0194[324] NET0194[325] NET0194[326] NET0194[327] 
+ NET0194[328] NET0194[329] NET0194[330] NET0194[331] NET0194[332] 
+ NET0194[333] NET0194[334] NET0194[335] NET0194[336] NET0194[337] 
+ NET0194[338] NET0194[339] NET0194[340] NET0194[341] NET0194[342] 
+ NET0194[343] NET0194[344] NET0194[345] NET0194[346] NET0194[347] 
+ NET0194[348] NET0194[349] NET0194[350] NET0194[351] NET0194[352] 
+ NET0194[353] NET0194[354] NET0194[355] NET0194[356] NET0194[357] 
+ NET0194[358] NET0194[359] NET0194[360] NET0194[361] NET0194[362] 
+ NET0194[363] NET0194[364] NET0194[365] NET0194[366] NET0194[367] 
+ NET0194[368] NET0194[369] NET0194[370] NET0194[371] NET0194[372] 
+ NET0194[373] NET0194[374] NET0194[375] NET0194[376] NET0194[377] 
+ NET0194[378] NET0194[379] NET0194[380] NET0194[381] NET0194[382] 
+ NET0194[383] NET0194[384] NET0194[385] NET0194[386] NET0194[387] 
+ NET0194[388] NET0194[389] NET0194[390] NET0194[391] NET0194[392] 
+ NET0194[393] NET0194[394] NET0194[395] NET0194[396] NET0194[397] 
+ NET0194[398] NET0194[399] NET0194[400] NET0194[401] NET0194[402] 
+ NET0194[403] NET0194[404] NET0194[405] NET0194[406] NET0194[407] 
+ NET0194[408] NET0194[409] NET0194[410] NET0194[411] NET0194[412] 
+ NET0194[413] NET0194[414] NET0194[415] NET0194[416] NET0194[417] 
+ NET0194[418] NET0194[419] NET0194[420] NET0194[421] NET0194[422] 
+ NET0194[423] NET0194[424] NET0194[425] NET0194[426] NET0194[427] 
+ NET0194[428] NET0194[429] NET0194[430] NET0194[431] NET0194[432] 
+ NET0194[433] NET0194[434] NET0194[435] NET0194[436] NET0194[437] 
+ NET0194[438] NET0194[439] NET0194[440] NET0194[441] NET0194[442] 
+ NET0194[443] NET0194[444] NET0194[445] NET0194[446] NET0194[447] 
+ NET0194[448] NET0194[449] NET0194[450] NET0194[451] NET0194[452] 
+ NET0194[453] NET0194[454] NET0194[455] NET0194[456] NET0194[457] 
+ NET0194[458] NET0194[459] NET0194[460] NET0194[461] NET0194[462] 
+ NET0194[463] NET0194[464] NET0194[465] NET0194[466] NET0194[467] 
+ NET0194[468] NET0194[469] NET0194[470] NET0194[471] NET0194[472] 
+ NET0194[473] NET0194[474] NET0194[475] NET0194[476] NET0194[477] 
+ NET0194[478] NET0194[479] NET0194[480] NET0194[481] NET0194[482] 
+ NET0194[483] NET0194[484] NET0194[485] NET0194[486] NET0194[487] 
+ NET0194[488] NET0194[489] NET0194[490] NET0194[491] NET0194[492] 
+ NET0194[493] NET0194[494] NET0194[495] NET0194[496] NET0194[497] 
+ NET0194[498] NET0194[499] NET0194[500] NET0194[501] NET0194[502] 
+ NET0194[503] NET0194[504] NET0194[505] NET0194[506] NET0194[507] 
+ NET0194[508] NET0194[509] NET0194[510] NET0194[511] NET01 NET21[0] NET21[1] 
+ NET21[2] NET14[0] NET14[1] NET14[2] NET14[3] NET14[4] NET14[5] NET14[6] 
+ NET14[7] NET14[8] NET13[0] NET13[1] NET13[2] NET13[3] NET13[4] NET13[5] 
+ NET13[6] NET13[7] NET13[8] NET4[0] NET4[1] NET4[2] NET4[3] NET3[0] NET3[1] 
+ NET3[2] NET3[3] S1AHSF400W40_SIM_SB
XI0 NET169 NET168 NET166 NET162 NET161 NET148 NET165 NET164 NET163 NET147 
+ NET146 NET145 NET144 NET176[0] NET176[1] NET176[2] NET176[3] NET176[4] 
+ NET176[5] NET176[6] NET176[7] NET176[8] NET176[9] NET176[10] NET175[0] 
+ NET175[1] NET175[2] NET175[3] NET175[4] NET175[5] NET175[6] NET175[7] 
+ NET175[8] NET175[9] NET175[10] NET159 NET158 NET172 NET171 NET157 NET156 
+ NET155 NET174[0] NET174[1] NET153 NET152 NET170 NET151 NET141 NET140 NET150 
+ NET149 NET0224[0] NET0224[1] NET0224[2] NET0224[3] NET0224[4] NET0224[5] 
+ NET0224[6] NET0224[7] NET0224[8] NET0224[9] NET0224[10] NET0224[11] 
+ NET0224[12] NET0224[13] NET0224[14] NET0224[15] NET0224[16] NET0224[17] 
+ NET0224[18] NET0224[19] NET0224[20] NET0224[21] NET0224[22] NET0224[23] 
+ NET0224[24] NET0224[25] NET0224[26] NET0224[27] NET0224[28] NET0224[29] 
+ NET0224[30] NET0224[31] NET0224[32] NET0224[33] NET0224[34] NET0224[35] 
+ NET0224[36] NET0224[37] NET0224[38] NET0224[39] NET0224[40] NET0224[41] 
+ NET0224[42] NET0224[43] NET0224[44] NET0224[45] NET0224[46] NET0224[47] 
+ NET0224[48] NET0224[49] NET0224[50] NET0224[51] NET0224[52] NET0224[53] 
+ NET0224[54] NET0224[55] NET0224[56] NET0224[57] NET0224[58] NET0224[59] 
+ NET0224[60] NET0224[61] NET0224[62] NET0224[63] NET0224[64] NET0224[65] 
+ NET0224[66] NET0224[67] NET0224[68] NET0224[69] NET0224[70] NET0224[71] 
+ NET0224[72] NET0224[73] NET0224[74] NET0224[75] NET0224[76] NET0224[77] 
+ NET0224[78] NET0224[79] NET0224[80] NET0224[81] NET0224[82] NET0224[83] 
+ NET0224[84] NET0224[85] NET0224[86] NET0224[87] NET0224[88] NET0224[89] 
+ NET0224[90] NET0224[91] NET0224[92] NET0224[93] NET0224[94] NET0224[95] 
+ NET0224[96] NET0224[97] NET0224[98] NET0224[99] NET0224[100] NET0224[101] 
+ NET0224[102] NET0224[103] NET0224[104] NET0224[105] NET0224[106] 
+ NET0224[107] NET0224[108] NET0224[109] NET0224[110] NET0224[111] 
+ NET0224[112] NET0224[113] NET0224[114] NET0224[115] NET0224[116] 
+ NET0224[117] NET0224[118] NET0224[119] NET0224[120] NET0224[121] 
+ NET0224[122] NET0224[123] NET0224[124] NET0224[125] NET0224[126] 
+ NET0224[127] NET0224[128] NET0224[129] NET0224[130] NET0224[131] 
+ NET0224[132] NET0224[133] NET0224[134] NET0224[135] NET0224[136] 
+ NET0224[137] NET0224[138] NET0224[139] NET0224[140] NET0224[141] 
+ NET0224[142] NET0224[143] NET0224[144] NET0224[145] NET0224[146] 
+ NET0224[147] NET0224[148] NET0224[149] NET0224[150] NET0224[151] 
+ NET0224[152] NET0224[153] NET0224[154] NET0224[155] NET0224[156] 
+ NET0224[157] NET0224[158] NET0224[159] NET0224[160] NET0224[161] 
+ NET0224[162] NET0224[163] NET0224[164] NET0224[165] NET0224[166] 
+ NET0224[167] NET0224[168] NET0224[169] NET0224[170] NET0224[171] 
+ NET0224[172] NET0224[173] NET0224[174] NET0224[175] NET0224[176] 
+ NET0224[177] NET0224[178] NET0224[179] NET0224[180] NET0224[181] 
+ NET0224[182] NET0224[183] NET0224[184] NET0224[185] NET0224[186] 
+ NET0224[187] NET0224[188] NET0224[189] NET0224[190] NET0224[191] 
+ NET0224[192] NET0224[193] NET0224[194] NET0224[195] NET0224[196] 
+ NET0224[197] NET0224[198] NET0224[199] NET0224[200] NET0224[201] 
+ NET0224[202] NET0224[203] NET0224[204] NET0224[205] NET0224[206] 
+ NET0224[207] NET0224[208] NET0224[209] NET0224[210] NET0224[211] 
+ NET0224[212] NET0224[213] NET0224[214] NET0224[215] NET0224[216] 
+ NET0224[217] NET0224[218] NET0224[219] NET0224[220] NET0224[221] 
+ NET0224[222] NET0224[223] NET0224[224] NET0224[225] NET0224[226] 
+ NET0224[227] NET0224[228] NET0224[229] NET0224[230] NET0224[231] 
+ NET0224[232] NET0224[233] NET0224[234] NET0224[235] NET0224[236] 
+ NET0224[237] NET0224[238] NET0224[239] NET0224[240] NET0224[241] 
+ NET0224[242] NET0224[243] NET0224[244] NET0224[245] NET0224[246] 
+ NET0224[247] NET0224[248] NET0224[249] NET0224[250] NET0224[251] 
+ NET0224[252] NET0224[253] NET0224[254] NET0224[255] NET0224[256] 
+ NET0224[257] NET0224[258] NET0224[259] NET0224[260] NET0224[261] 
+ NET0224[262] NET0224[263] NET0224[264] NET0224[265] NET0224[266] 
+ NET0224[267] NET0224[268] NET0224[269] NET0224[270] NET0224[271] 
+ NET0224[272] NET0224[273] NET0224[274] NET0224[275] NET0224[276] 
+ NET0224[277] NET0224[278] NET0224[279] NET0224[280] NET0224[281] 
+ NET0224[282] NET0224[283] NET0224[284] NET0224[285] NET0224[286] 
+ NET0224[287] NET0224[288] NET0224[289] NET0224[290] NET0224[291] 
+ NET0224[292] NET0224[293] NET0224[294] NET0224[295] NET0224[296] 
+ NET0224[297] NET0224[298] NET0224[299] NET0224[300] NET0224[301] 
+ NET0224[302] NET0224[303] NET0224[304] NET0224[305] NET0224[306] 
+ NET0224[307] NET0224[308] NET0224[309] NET0224[310] NET0224[311] 
+ NET0224[312] NET0224[313] NET0224[314] NET0224[315] NET0224[316] 
+ NET0224[317] NET0224[318] NET0224[319] NET0224[320] NET0224[321] 
+ NET0224[322] NET0224[323] NET0224[324] NET0224[325] NET0224[326] 
+ NET0224[327] NET0224[328] NET0224[329] NET0224[330] NET0224[331] 
+ NET0224[332] NET0224[333] NET0224[334] NET0224[335] NET0224[336] 
+ NET0224[337] NET0224[338] NET0224[339] NET0224[340] NET0224[341] 
+ NET0224[342] NET0224[343] NET0224[344] NET0224[345] NET0224[346] 
+ NET0224[347] NET0224[348] NET0224[349] NET0224[350] NET0224[351] 
+ NET0224[352] NET0224[353] NET0224[354] NET0224[355] NET0224[356] 
+ NET0224[357] NET0224[358] NET0224[359] NET0224[360] NET0224[361] 
+ NET0224[362] NET0224[363] NET0224[364] NET0224[365] NET0224[366] 
+ NET0224[367] NET0224[368] NET0224[369] NET0224[370] NET0224[371] 
+ NET0224[372] NET0224[373] NET0224[374] NET0224[375] NET0224[376] 
+ NET0224[377] NET0224[378] NET0224[379] NET0224[380] NET0224[381] 
+ NET0224[382] NET0224[383] NET0224[384] NET0224[385] NET0224[386] 
+ NET0224[387] NET0224[388] NET0224[389] NET0224[390] NET0224[391] 
+ NET0224[392] NET0224[393] NET0224[394] NET0224[395] NET0224[396] 
+ NET0224[397] NET0224[398] NET0224[399] NET0224[400] NET0224[401] 
+ NET0224[402] NET0224[403] NET0224[404] NET0224[405] NET0224[406] 
+ NET0224[407] NET0224[408] NET0224[409] NET0224[410] NET0224[411] 
+ NET0224[412] NET0224[413] NET0224[414] NET0224[415] NET0224[416] 
+ NET0224[417] NET0224[418] NET0224[419] NET0224[420] NET0224[421] 
+ NET0224[422] NET0224[423] NET0224[424] NET0224[425] NET0224[426] 
+ NET0224[427] NET0224[428] NET0224[429] NET0224[430] NET0224[431] 
+ NET0224[432] NET0224[433] NET0224[434] NET0224[435] NET0224[436] 
+ NET0224[437] NET0224[438] NET0224[439] NET0224[440] NET0224[441] 
+ NET0224[442] NET0224[443] NET0224[444] NET0224[445] NET0224[446] 
+ NET0224[447] NET0224[448] NET0224[449] NET0224[450] NET0224[451] 
+ NET0224[452] NET0224[453] NET0224[454] NET0224[455] NET0224[456] 
+ NET0224[457] NET0224[458] NET0224[459] NET0224[460] NET0224[461] 
+ NET0224[462] NET0224[463] NET0224[464] NET0224[465] NET0224[466] 
+ NET0224[467] NET0224[468] NET0224[469] NET0224[470] NET0224[471] 
+ NET0224[472] NET0224[473] NET0224[474] NET0224[475] NET0224[476] 
+ NET0224[477] NET0224[478] NET0224[479] NET0224[480] NET0224[481] 
+ NET0224[482] NET0224[483] NET0224[484] NET0224[485] NET0224[486] 
+ NET0224[487] NET0224[488] NET0224[489] NET0224[490] NET0224[491] 
+ NET0224[492] NET0224[493] NET0224[494] NET0224[495] NET0224[496] 
+ NET0224[497] NET0224[498] NET0224[499] NET0224[500] NET0224[501] 
+ NET0224[502] NET0224[503] NET0224[504] NET0224[505] NET0224[506] 
+ NET0224[507] NET0224[508] NET0224[509] NET0224[510] NET0224[511] NET031 
+ NET167[0] NET167[1] NET167[2] NET160[0] NET160[1] NET160[2] NET160[3] 
+ NET160[4] NET160[5] NET160[6] NET160[7] NET160[8] NET160[9] NET160[10] 
+ NET154[0] NET154[1] NET154[2] NET154[3] NET154[4] NET154[5] NET154[6] 
+ NET154[7] NET154[8] NET154[9] NET154[10] NET143[0] NET143[1] NET143[2] 
+ NET143[3] NET142[0] NET142[1] NET142[2] NET142[3] S1AHSF400W40_SIM_FULL
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MCNTIOX8_F
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCNTIOX8_F AWT BIST BLTRKWLDRV BWEB[0] BWEB[1] BWEB[2] BWEB[3] BWEB[4] 
+ BWEB[5] BWEB[6] BWEB[7] BWEBM[0] BWEBM[1] BWEBM[2] BWEBM[3] BWEBM[4] 
+ BWEBM[5] BWEBM[6] BWEBM[7] CEB CEBM CLK D[0] D[1] D[2] D[3] D[4] D[5] D[6] 
+ D[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] 
+ DM[0] DM[1] DM[2] DM[3] DM[4] DM[5] DM[6] DM[7] GBL[0] GBL[1] GBL[2] GBL[3] 
+ GBL[4] GBL[5] GBL[6] GBL[7] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] 
+ GBLB[6] GBLB[7] GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GWB[0] 
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] PD_BUF PD_CVDDBUF Q[0] Q[1] 
+ Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] REDEN REDENB RTSEL[0] RTSEL[1] RW_RE SLP TM 
+ TRKBL VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAE_TK WTSEL[0] WTSEL[1] 
+ WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] 
+ XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] 
+ YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I BWEB[0]:I BWEB[1]:I BWEB[2]:I BWEB[3]:I BWEB[4]:I 
*.PININFO BWEB[5]:I BWEB[6]:I BWEB[7]:I BWEBM[0]:I BWEBM[1]:I BWEBM[2]:I 
*.PININFO BWEBM[3]:I BWEBM[4]:I BWEBM[5]:I BWEBM[6]:I BWEBM[7]:I CEB:I CEBM:I 
*.PININFO CLK:I D[0]:I D[1]:I D[2]:I D[3]:I D[4]:I D[5]:I D[6]:I D[7]:I 
*.PININFO DM[0]:I DM[1]:I DM[2]:I DM[3]:I DM[4]:I DM[5]:I DM[6]:I DM[7]:I 
*.PININFO REDEN:I REDENB:I RTSEL[0]:I RTSEL[1]:I SLP:I TM:I WEB:I WEBM:I 
*.PININFO WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I 
*.PININFO X[5]:I X[6]:I X[7]:I X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I 
*.PININFO XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I 
*.PININFO Y[0]:I Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I Q[0]:O 
*.PININFO Q[1]:O Q[2]:O Q[3]:O Q[4]:O Q[5]:O Q[6]:O Q[7]:O VHI:O VLO:O 
*.PININFO BLTRKWLDRV:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B GBL[0]:B GBL[1]:B GBL[2]:B GBL[3]:B GBL[4]:B GBL[5]:B 
*.PININFO GBL[6]:B GBL[7]:B GBLB[0]:B GBLB[1]:B GBLB[2]:B GBLB[3]:B GBLB[4]:B 
*.PININFO GBLB[5]:B GBLB[6]:B GBLB[7]:B GW[0]:B GW[1]:B GW[2]:B GW[3]:B 
*.PININFO GW[4]:B GW[5]:B GW[6]:B GW[7]:B GWB[0]:B GWB[1]:B GWB[2]:B GWB[3]:B 
*.PININFO GWB[4]:B GWB[5]:B GWB[6]:B GWB[7]:B PD_BUF:B PD_CVDDBUF:B RW_RE:B 
*.PININFO TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XI8 AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] 
+ DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] SLP PD_BUF PD_CVDDBUF NET153 
+ REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL VDDHD VDDI VHI VLO VSSI WEB 
+ WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] 
+ X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] 
+ YM[3] S1AHSF400W40_CNT_CORE_F_M4
XIO_M8_L<0> AWT2 BIST2IO BWEB[0] BWEBM[0] CKD D[0] DM[0] GBL[0] GBLB[0] GW[0] 
+ GWB[0] PD_BUF Q[0] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XIO_M8_L<1> AWT2 BIST2IO BWEB[1] BWEBM[1] CKD D[1] DM[1] GBL[1] GBLB[1] GW[1] 
+ GWB[1] PD_BUF Q[1] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XIO_M8_L<2> AWT2 BIST2IO BWEB[2] BWEBM[2] CKD D[2] DM[2] GBL[2] GBLB[2] GW[2] 
+ GWB[2] PD_BUF Q[2] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XIO_M8_L<3> AWT2 BIST2IO BWEB[3] BWEBM[3] CKD D[3] DM[3] GBL[3] GBLB[3] GW[3] 
+ GWB[3] PD_BUF Q[3] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XI2<4> AWT2 BIST2IO BWEB[4] BWEBM[4] CKD D[4] DM[4] GBL[4] GBLB[4] GW[4] 
+ GWB[4] PD_BUF Q[4] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XI2<5> AWT2 BIST2IO BWEB[5] BWEBM[5] CKD D[5] DM[5] GBL[5] GBLB[5] GW[5] 
+ GWB[5] PD_BUF Q[5] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XI2<6> AWT2 BIST2IO BWEB[6] BWEBM[6] CKD D[6] DM[6] GBL[6] GBLB[6] GW[6] 
+ GWB[6] PD_BUF Q[6] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XI2<7> AWT2 BIST2IO BWEB[7] BWEBM[7] CKD D[7] DM[7] GBL[7] GBLB[7] GW[7] 
+ GWB[7] PD_BUF Q[7] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MCNTIOX2_F
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCNTIOX2_F AWT BIST BLTRKWLDRV BWEB[0] BWEB[1] BWEBM[0] BWEBM[1] CEB 
+ CEBM CLK D[0] D[1] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] 
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DM[0] DM[1] GBL[0] GBL[1] GBLB[0] GBLB[1] GW[0] GW[1] 
+ GWB[0] GWB[1] PD_BUF PD_CVDDBUF Q[0] Q[1] REDEN REDENB RTSEL[0] RTSEL[1] 
+ RW_RE SLP TM TRKBL VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] 
+ X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] 
+ Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I BWEB[0]:I BWEB[1]:I BWEBM[0]:I BWEBM[1]:I CEB:I CEBM:I 
*.PININFO CLK:I D[0]:I D[1]:I DM[0]:I DM[1]:I REDEN:I REDENB:I RTSEL[0]:I 
*.PININFO RTSEL[1]:I SLP:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I 
*.PININFO X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I 
*.PININFO X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I XM[5]:I 
*.PININFO XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I Y[2]:I Y[3]:I 
*.PININFO YM[0]:I YM[1]:I YM[2]:I YM[3]:I Q[0]:O Q[1]:O VHI:O VLO:O 
*.PININFO BLTRKWLDRV:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B GBL[0]:B GBL[1]:B GBLB[0]:B GBLB[1]:B GW[0]:B GW[1]:B 
*.PININFO GWB[0]:B GWB[1]:B PD_BUF:B PD_CVDDBUF:B RW_RE:B TRKBL:B VDDHD:B 
*.PININFO VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XI0 AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] 
+ DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] SLP PD_BUF PD_CVDDBUF NET86 
+ REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL VDDHD VDDI VHI VLO VSSI WEB 
+ WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] 
+ X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] 
+ YM[3] S1AHSF400W40_CNT_CORE_F_M16
XIO_M4_L AWT2 BIST2IO BWEB[0] BWEBM[0] CKD D[0] DM[0] GBL[0] GBLB[0] GW[0] 
+ GWB[0] PD_BUF Q[0] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M16
XI2 AWT2 BIST2IO BWEB[1] BWEBM[1] CKD D[1] DM[1] GBL[1] GBLB[1] GW[1] GWB[1] 
+ PD_BUF Q[1] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M16
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MCNTIOX4_F
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCNTIOX4_F AWT BIST BLTRKWLDRV BWEB[0] BWEB[1] BWEB[2] BWEB[3] 
+ BWEBM[0] BWEBM[1] BWEBM[2] BWEBM[3] CEB CEBM CLK D[0] D[1] D[2] D[3] 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] 
+ DM[0] DM[1] DM[2] DM[3] GBL[0] GBL[1] GBL[2] GBL[3] GBLB[0] GBLB[1] GBLB[2] 
+ GBLB[3] GW[0] GW[1] GW[2] GW[3] GWB[0] GWB[1] GWB[2] GWB[3] PD_BUF 
+ PD_CVDDBUF Q[0] Q[1] Q[2] Q[3] REDEN REDENB RTSEL[0] RTSEL[1] RW_RE SLP TM 
+ TRKBL VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAE_TK WTSEL[0] WTSEL[1] 
+ WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] 
+ XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] 
+ YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I BWEB[0]:I BWEB[1]:I BWEB[2]:I BWEB[3]:I BWEBM[0]:I 
*.PININFO BWEBM[1]:I BWEBM[2]:I BWEBM[3]:I CEB:I CEBM:I CLK:I D[0]:I D[1]:I 
*.PININFO D[2]:I D[3]:I DM[0]:I DM[1]:I DM[2]:I DM[3]:I REDEN:I REDENB:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I SLP:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I 
*.PININFO XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I 
*.PININFO Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I Q[0]:O Q[1]:O Q[2]:O 
*.PININFO Q[3]:O VHI:O VLO:O BLTRKWLDRV:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B 
*.PININFO DEC_X0[3]:B DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B 
*.PININFO DEC_X1[0]:B DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B 
*.PININFO DEC_X1[5]:B DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B 
*.PININFO DEC_X2[2]:B DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B 
*.PININFO DEC_X3[3]:B DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B 
*.PININFO DEC_Y[0]:B DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B 
*.PININFO DEC_Y[6]:B DEC_Y[7]:B GBL[0]:B GBL[1]:B GBL[2]:B GBL[3]:B GBLB[0]:B 
*.PININFO GBLB[1]:B GBLB[2]:B GBLB[3]:B GW[0]:B GW[1]:B GW[2]:B GW[3]:B 
*.PININFO GWB[0]:B GWB[1]:B GWB[2]:B GWB[3]:B PD_BUF:B PD_CVDDBUF:B RW_RE:B 
*.PININFO TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XI7 AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] 
+ DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] SLP PD_BUF PD_CVDDBUF NET86 
+ REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL VDDHD VDDI VHI VLO VSSI WEB 
+ WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] 
+ X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] 
+ YM[3] S1AHSF400W40_CNT_CORE_F_M8
XIO_M8_L<0> AWT2 BIST2IO BWEB[0] BWEBM[0] CKD D[0] DM[0] GBL[0] GBLB[0] GW[0] 
+ GWB[0] PD_BUF Q[0] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M8
XIO_M8_L<1> AWT2 BIST2IO BWEB[1] BWEBM[1] CKD D[1] DM[1] GBL[1] GBLB[1] GW[1] 
+ GWB[1] PD_BUF Q[1] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M8
XI2<2> AWT2 BIST2IO BWEB[2] BWEBM[2] CKD D[2] DM[2] GBL[2] GBLB[2] GW[2] 
+ GWB[2] PD_BUF Q[2] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M8
XI2<3> AWT2 BIST2IO BWEB[3] BWEBM[3] CKD D[3] DM[3] GBL[3] GBLB[3] GW[3] 
+ GWB[3] PD_BUF Q[3] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M8
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MCNTIOX2_F_BIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCNTIOX2_F_BIST AWT BIST BLTRKWLDRV BWEB[0] BWEB[1] BWEBM[0] BWEBM[1] 
+ CEB CEBM CLK D[0] D[1] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] 
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DM[0] DM[1] GBL[0] GBL[1] GBLB[0] GBLB[1] GW[0] GW[1] 
+ GWB[0] GWB[1] PD_BUF PD_CVDDBUF Q[0] Q[1] REDEN REDENB RTSEL[0] RTSEL[1] 
+ RW_RE SLP TM TRKBL VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] 
+ X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] 
+ Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I BWEB[0]:I BWEB[1]:I BWEBM[0]:I BWEBM[1]:I CEB:I CEBM:I 
*.PININFO CLK:I D[0]:I D[1]:I DM[0]:I DM[1]:I REDEN:I REDENB:I RTSEL[0]:I 
*.PININFO RTSEL[1]:I SLP:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I 
*.PININFO X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I 
*.PININFO X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I XM[5]:I 
*.PININFO XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I Y[2]:I Y[3]:I 
*.PININFO YM[0]:I YM[1]:I YM[2]:I YM[3]:I Q[0]:O Q[1]:O VHI:O VLO:O 
*.PININFO BLTRKWLDRV:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B GBL[0]:B GBL[1]:B GBLB[0]:B GBLB[1]:B GW[0]:B GW[1]:B 
*.PININFO GWB[0]:B GWB[1]:B PD_BUF:B PD_CVDDBUF:B RW_RE:B TRKBL:B VDDHD:B 
*.PININFO VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XI0 AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] 
+ DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] SLP PD_BUF PD_CVDDBUF NET86 
+ REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL VDDHD VDDI VHI VLO VSSI WEB 
+ WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] 
+ X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] 
+ YM[3] S1AHSF400W40_CNT_CORE_F_M16_BIST
XIO_M4_L AWT2 BIST2IO BWEB[0] BWEBM[0] CKD D[0] DM[0] GBL[0] GBLB[0] GW[0] 
+ GWB[0] PD_BUF Q[0] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M16
XI2 AWT2 BIST2IO BWEB[1] BWEBM[1] CKD D[1] DM[1] GBL[1] GBLB[1] GW[1] GWB[1] 
+ PD_BUF Q[1] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M16
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MCNTIOX4_F_BIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCNTIOX4_F_BIST AWT BIST BLTRKWLDRV BWEB[0] BWEB[1] BWEB[2] BWEB[3] 
+ BWEBM[0] BWEBM[1] BWEBM[2] BWEBM[3] CEB CEBM CLK D[0] D[1] D[2] D[3] 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] 
+ DM[0] DM[1] DM[2] DM[3] GBL[0] GBL[1] GBL[2] GBL[3] GBLB[0] GBLB[1] GBLB[2] 
+ GBLB[3] GW[0] GW[1] GW[2] GW[3] GWB[0] GWB[1] GWB[2] GWB[3] PD_BUF 
+ PD_CVDDBUF Q[0] Q[1] Q[2] Q[3] REDEN REDENB RTSEL[0] RTSEL[1] RW_RE SLP TM 
+ TRKBL VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAE_TK WTSEL[0] WTSEL[1] 
+ WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] 
+ XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] 
+ YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I BWEB[0]:I BWEB[1]:I BWEB[2]:I BWEB[3]:I BWEBM[0]:I 
*.PININFO BWEBM[1]:I BWEBM[2]:I BWEBM[3]:I CEB:I CEBM:I CLK:I D[0]:I D[1]:I 
*.PININFO D[2]:I D[3]:I DM[0]:I DM[1]:I DM[2]:I DM[3]:I REDEN:I REDENB:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I SLP:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I 
*.PININFO XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I 
*.PININFO Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I Q[0]:O Q[1]:O Q[2]:O 
*.PININFO Q[3]:O VHI:O VLO:O BLTRKWLDRV:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B 
*.PININFO DEC_X0[3]:B DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B 
*.PININFO DEC_X1[0]:B DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B 
*.PININFO DEC_X1[5]:B DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B 
*.PININFO DEC_X2[2]:B DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B 
*.PININFO DEC_X3[3]:B DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B 
*.PININFO DEC_Y[0]:B DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B 
*.PININFO DEC_Y[6]:B DEC_Y[7]:B GBL[0]:B GBL[1]:B GBL[2]:B GBL[3]:B GBLB[0]:B 
*.PININFO GBLB[1]:B GBLB[2]:B GBLB[3]:B GW[0]:B GW[1]:B GW[2]:B GW[3]:B 
*.PININFO GWB[0]:B GWB[1]:B GWB[2]:B GWB[3]:B PD_BUF:B PD_CVDDBUF:B RW_RE:B 
*.PININFO TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XI7 AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] 
+ DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] SLP PD_BUF PD_CVDDBUF NET86 
+ REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL VDDHD VDDI VHI VLO VSSI WEB 
+ WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] 
+ X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] 
+ YM[3] S1AHSF400W40_CNT_CORE_F_M8_BIST
XIO_M8_L<0> AWT2 BIST2IO BWEB[0] BWEBM[0] CKD D[0] DM[0] GBL[0] GBLB[0] GW[0] 
+ GWB[0] PD_BUF Q[0] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M8
XIO_M8_L<1> AWT2 BIST2IO BWEB[1] BWEBM[1] CKD D[1] DM[1] GBL[1] GBLB[1] GW[1] 
+ GWB[1] PD_BUF Q[1] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M8
XI2<2> AWT2 BIST2IO BWEB[2] BWEBM[2] CKD D[2] DM[2] GBL[2] GBLB[2] GW[2] 
+ GWB[2] PD_BUF Q[2] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M8
XI2<3> AWT2 BIST2IO BWEB[3] BWEBM[3] CKD D[3] DM[3] GBL[3] GBLB[3] GW[3] 
+ GWB[3] PD_BUF Q[3] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M8
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MCNTIOX8_F_BIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCNTIOX8_F_BIST AWT BIST BLTRKWLDRV BWEB[0] BWEB[1] BWEB[2] BWEB[3] 
+ BWEB[4] BWEB[5] BWEB[6] BWEB[7] BWEBM[0] BWEBM[1] BWEBM[2] BWEBM[3] BWEBM[4] 
+ BWEBM[5] BWEBM[6] BWEBM[7] CEB CEBM CLK D[0] D[1] D[2] D[3] D[4] D[5] D[6] 
+ D[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] 
+ DM[0] DM[1] DM[2] DM[3] DM[4] DM[5] DM[6] DM[7] GBL[0] GBL[1] GBL[2] GBL[3] 
+ GBL[4] GBL[5] GBL[6] GBL[7] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] 
+ GBLB[6] GBLB[7] GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GWB[0] 
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] PD_BUF PD_CVDDBUF Q[0] Q[1] 
+ Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] REDEN REDENB RTSEL[0] RTSEL[1] RW_RE SLP TM 
+ TRKBL VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAE_TK WTSEL[0] WTSEL[1] 
+ WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] 
+ XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] 
+ YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I BWEB[0]:I BWEB[1]:I BWEB[2]:I BWEB[3]:I BWEB[4]:I 
*.PININFO BWEB[5]:I BWEB[6]:I BWEB[7]:I BWEBM[0]:I BWEBM[1]:I BWEBM[2]:I 
*.PININFO BWEBM[3]:I BWEBM[4]:I BWEBM[5]:I BWEBM[6]:I BWEBM[7]:I CEB:I CEBM:I 
*.PININFO CLK:I D[0]:I D[1]:I D[2]:I D[3]:I D[4]:I D[5]:I D[6]:I D[7]:I 
*.PININFO DM[0]:I DM[1]:I DM[2]:I DM[3]:I DM[4]:I DM[5]:I DM[6]:I DM[7]:I 
*.PININFO REDEN:I REDENB:I RTSEL[0]:I RTSEL[1]:I SLP:I TM:I WEB:I WEBM:I 
*.PININFO WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I 
*.PININFO X[5]:I X[6]:I X[7]:I X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I 
*.PININFO XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I 
*.PININFO Y[0]:I Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I Q[0]:O 
*.PININFO Q[1]:O Q[2]:O Q[3]:O Q[4]:O Q[5]:O Q[6]:O Q[7]:O VHI:O VLO:O 
*.PININFO BLTRKWLDRV:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B GBL[0]:B GBL[1]:B GBL[2]:B GBL[3]:B GBL[4]:B GBL[5]:B 
*.PININFO GBL[6]:B GBL[7]:B GBLB[0]:B GBLB[1]:B GBLB[2]:B GBLB[3]:B GBLB[4]:B 
*.PININFO GBLB[5]:B GBLB[6]:B GBLB[7]:B GW[0]:B GW[1]:B GW[2]:B GW[3]:B 
*.PININFO GW[4]:B GW[5]:B GW[6]:B GW[7]:B GWB[0]:B GWB[1]:B GWB[2]:B GWB[3]:B 
*.PININFO GWB[4]:B GWB[5]:B GWB[6]:B GWB[7]:B PD_BUF:B PD_CVDDBUF:B RW_RE:B 
*.PININFO TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XI8 AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] 
+ DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] SLP PD_BUF PD_CVDDBUF NET153 
+ REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL VDDHD VDDI VHI VLO VSSI WEB 
+ WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] 
+ X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] 
+ YM[3] S1AHSF400W40_CNT_CORE_F_M4_BIST
XIO_M8_L<0> AWT2 BIST2IO BWEB[0] BWEBM[0] CKD D[0] DM[0] GBL[0] GBLB[0] GW[0] 
+ GWB[0] PD_BUF Q[0] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XIO_M8_L<1> AWT2 BIST2IO BWEB[1] BWEBM[1] CKD D[1] DM[1] GBL[1] GBLB[1] GW[1] 
+ GWB[1] PD_BUF Q[1] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XIO_M8_L<2> AWT2 BIST2IO BWEB[2] BWEBM[2] CKD D[2] DM[2] GBL[2] GBLB[2] GW[2] 
+ GWB[2] PD_BUF Q[2] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XIO_M8_L<3> AWT2 BIST2IO BWEB[3] BWEBM[3] CKD D[3] DM[3] GBL[3] GBLB[3] GW[3] 
+ GWB[3] PD_BUF Q[3] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XI2<4> AWT2 BIST2IO BWEB[4] BWEBM[4] CKD D[4] DM[4] GBL[4] GBLB[4] GW[4] 
+ GWB[4] PD_BUF Q[4] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XI2<5> AWT2 BIST2IO BWEB[5] BWEBM[5] CKD D[5] DM[5] GBL[5] GBLB[5] GW[5] 
+ GWB[5] PD_BUF Q[5] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XI2<6> AWT2 BIST2IO BWEB[6] BWEBM[6] CKD D[6] DM[6] GBL[6] GBLB[6] GW[6] 
+ GWB[6] PD_BUF Q[6] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XI2<7> AWT2 BIST2IO BWEB[7] BWEBM[7] CKD D[7] DM[7] GBL[7] GBLB[7] GW[7] 
+ GWB[7] PD_BUF Q[7] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    MCB_2X16_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_2X16_CHAR BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] 
+ BL[9] BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BLB[0] BLB[1] BLB[2] BLB[3] 
+ BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] 
+ BLB[14] BLB[15] GBL GBLB GW GWB VDDI VSSI WL[0] WL[1]
*.PININFO WL[0]:I WL[1]:I BL[0]:B BL[1]:B BL[2]:B BL[3]:B BL[4]:B BL[5]:B 
*.PININFO BL[6]:B BL[7]:B BL[8]:B BL[9]:B BL[10]:B BL[11]:B BL[12]:B BL[13]:B 
*.PININFO BL[14]:B BL[15]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B BLB[4]:B 
*.PININFO BLB[5]:B BLB[6]:B BLB[7]:B BLB[8]:B BLB[9]:B BLB[10]:B BLB[11]:B 
*.PININFO BLB[12]:B BLB[13]:B BLB[14]:B BLB[15]:B GBL:B GBLB:B GW:B GWB:B 
*.PININFO VDDI:B VSSI:B
XMCB_1<0> BL[0] BLB[0] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<1> BL[1] BLB[1] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<2> BL[2] BLB[2] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<3> BL[3] BLB[3] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<4> BL[4] BLB[4] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<5> BL[5] BLB[5] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<6> BL[6] BLB[6] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<7> BL[7] BLB[7] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<8> BL[8] BLB[8] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<9> BL[9] BLB[9] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<10> BL[10] BLB[10] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<11> BL[11] BLB[11] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<12> BL[12] BLB[12] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<13> BL[13] BLB[13] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<14> BL[14] BLB[14] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<15> BL[15] BLB[15] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_0<0> BL[0] BLB[0] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<1> BL[1] BLB[1] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<2> BL[2] BLB[2] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<3> BL[3] BLB[3] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<4> BL[4] BLB[4] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<5> BL[5] BLB[5] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<6> BL[6] BLB[6] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<7> BL[7] BLB[7] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<8> BL[8] BLB[8] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<9> BL[9] BLB[9] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<10> BL[10] BLB[10] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<11> BL[11] BLB[11] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<12> BL[12] BLB[12] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<13> BL[13] BLB[13] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<14> BL[14] BLB[14] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<15> BL[15] BLB[15] VDDI VSSI WL[0] S1AHSF400W40_MCB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_CHAR
* CELL NAME:    MCB_2X8_CHAR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_2X8_CHAR BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BLB[0] 
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] GBL GBLB GW GWB VDDI VSSI 
+ WL[0] WL[1]
*.PININFO WL[0]:I WL[1]:I BL[0]:B BL[1]:B BL[2]:B BL[3]:B BL[4]:B BL[5]:B 
*.PININFO BL[6]:B BL[7]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B BLB[4]:B 
*.PININFO BLB[5]:B BLB[6]:B BLB[7]:B GBL:B GBLB:B GW:B GWB:B VDDI:B VSSI:B
XMCB_0<0> BL[0] BLB[0] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<1> BL[1] BLB[1] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<2> BL[2] BLB[2] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<3> BL[3] BLB[3] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<4> BL[4] BLB[4] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<5> BL[5] BLB[5] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<6> BL[6] BLB[6] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<7> BL[7] BLB[7] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_1<0> BL[0] BLB[0] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<1> BL[1] BLB[1] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<2> BL[2] BLB[2] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<3> BL[3] BLB[3] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<4> BL[4] BLB[4] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<5> BL[5] BLB[5] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<6> BL[6] BLB[6] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<7> BL[7] BLB[7] VDDI VSSI WL[1] S1AHSF400W40_MCB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MCB_2X16_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_2X16_SB BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] 
+ BL[9] BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BLB[0] BLB[1] BLB[2] BLB[3] 
+ BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] 
+ BLB[14] BLB[15] VDDI VSSI WL[0] WL[1]
*.PININFO WL[0]:I WL[1]:I BL[0]:B BL[1]:B BL[2]:B BL[3]:B BL[4]:B BL[5]:B 
*.PININFO BL[6]:B BL[7]:B BL[8]:B BL[9]:B BL[10]:B BL[11]:B BL[12]:B BL[13]:B 
*.PININFO BL[14]:B BL[15]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B BLB[4]:B 
*.PININFO BLB[5]:B BLB[6]:B BLB[7]:B BLB[8]:B BLB[9]:B BLB[10]:B BLB[11]:B 
*.PININFO BLB[12]:B BLB[13]:B BLB[14]:B BLB[15]:B VDDI:B VSSI:B
XMCB_1<0> BL[0] BLB[0] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<1> BL[1] BLB[1] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<2> BL[2] BLB[2] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<3> BL[3] BLB[3] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<4> BL[4] BLB[4] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<5> BL[5] BLB[5] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<6> BL[6] BLB[6] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<7> BL[7] BLB[7] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<8> BL[8] BLB[8] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<9> BL[9] BLB[9] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<10> BL[10] BLB[10] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<11> BL[11] BLB[11] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<12> BL[12] BLB[12] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<13> BL[13] BLB[13] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<14> BL[14] BLB[14] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<15> BL[15] BLB[15] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_0<0> BL[0] BLB[0] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<1> BL[1] BLB[1] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<2> BL[2] BLB[2] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<3> BL[3] BLB[3] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<4> BL[4] BLB[4] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<5> BL[5] BLB[5] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<6> BL[6] BLB[6] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<7> BL[7] BLB[7] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<8> BL[8] BLB[8] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<9> BL[9] BLB[9] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<10> BL[10] BLB[10] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<11> BL[11] BLB[11] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<12> BL[12] BLB[12] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<13> BL[13] BLB[13] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<14> BL[14] BLB[14] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<15> BL[15] BLB[15] VDDI VSSI WL[0] S1AHSF400W40_MCB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MCB_2X8_SB
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_2X8_SB BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BLB[0] 
+ BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] VDDI VSSI WL[0] WL[1]
*.PININFO WL[0]:I WL[1]:I BL[0]:B BL[1]:B BL[2]:B BL[3]:B BL[4]:B BL[5]:B 
*.PININFO BL[6]:B BL[7]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B BLB[4]:B 
*.PININFO BLB[5]:B BLB[6]:B BLB[7]:B VDDI:B VSSI:B
XMCB_0<0> BL[0] BLB[0] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<1> BL[1] BLB[1] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<2> BL[2] BLB[2] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<3> BL[3] BLB[3] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<4> BL[4] BLB[4] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<5> BL[5] BLB[5] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<6> BL[6] BLB[6] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<7> BL[7] BLB[7] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_1<0> BL[0] BLB[0] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<1> BL[1] BLB[1] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<2> BL[2] BLB[2] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<3> BL[3] BLB[3] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<4> BL[4] BLB[4] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<5> BL[5] BLB[5] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<6> BL[6] BLB[6] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<7> BL[7] BLB[7] VDDI VSSI WL[1] S1AHSF400W40_MCB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MCB_2X16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_2X16 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] 
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] 
+ BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] 
+ BLB[15] GBL GBLB GW GWB VDDI VSSI WL[0] WL[1]
*.PININFO WL[0]:I WL[1]:I BL[0]:B BL[1]:B BL[2]:B BL[3]:B BL[4]:B BL[5]:B 
*.PININFO BL[6]:B BL[7]:B BL[8]:B BL[9]:B BL[10]:B BL[11]:B BL[12]:B BL[13]:B 
*.PININFO BL[14]:B BL[15]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B BLB[4]:B 
*.PININFO BLB[5]:B BLB[6]:B BLB[7]:B BLB[8]:B BLB[9]:B BLB[10]:B BLB[11]:B 
*.PININFO BLB[12]:B BLB[13]:B BLB[14]:B BLB[15]:B GBL:B GBLB:B GW:B GWB:B 
*.PININFO VDDI:B VSSI:B
XMCB_1<0> BL[0] BLB[0] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<1> BL[1] BLB[1] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<2> BL[2] BLB[2] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<3> BL[3] BLB[3] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<4> BL[4] BLB[4] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<5> BL[5] BLB[5] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<6> BL[6] BLB[6] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<7> BL[7] BLB[7] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<8> BL[8] BLB[8] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<9> BL[9] BLB[9] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<10> BL[10] BLB[10] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<11> BL[11] BLB[11] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<12> BL[12] BLB[12] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<13> BL[13] BLB[13] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<14> BL[14] BLB[14] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<15> BL[15] BLB[15] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_0<0> BL[0] BLB[0] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<1> BL[1] BLB[1] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<2> BL[2] BLB[2] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<3> BL[3] BLB[3] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<4> BL[4] BLB[4] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<5> BL[5] BLB[5] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<6> BL[6] BLB[6] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<7> BL[7] BLB[7] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<8> BL[8] BLB[8] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<9> BL[9] BLB[9] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<10> BL[10] BLB[10] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<11> BL[11] BLB[11] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<12> BL[12] BLB[12] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<13> BL[13] BLB[13] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<14> BL[14] BLB[14] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<15> BL[15] BLB[15] VDDI VSSI WL[0] S1AHSF400W40_MCB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MCB_2X8
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_2X8 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BLB[0] BLB[1] 
+ BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] GBL GBLB GW GWB VDDI VSSI WL[0] 
+ WL[1]
*.PININFO WL[0]:I WL[1]:I BL[0]:B BL[1]:B BL[2]:B BL[3]:B BL[4]:B BL[5]:B 
*.PININFO BL[6]:B BL[7]:B BLB[0]:B BLB[1]:B BLB[2]:B BLB[3]:B BLB[4]:B 
*.PININFO BLB[5]:B BLB[6]:B BLB[7]:B GBL:B GBLB:B GW:B GWB:B VDDI:B VSSI:B
XMCB_0<0> BL[0] BLB[0] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<1> BL[1] BLB[1] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<2> BL[2] BLB[2] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<3> BL[3] BLB[3] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<4> BL[4] BLB[4] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<5> BL[5] BLB[5] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<6> BL[6] BLB[6] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_0<7> BL[7] BLB[7] VDDI VSSI WL[0] S1AHSF400W40_MCB
XMCB_1<0> BL[0] BLB[0] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<1> BL[1] BLB[1] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<2> BL[2] BLB[2] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<3> BL[3] BLB[3] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<4> BL[4] BLB[4] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<5> BL[5] BLB[5] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<6> BL[6] BLB[6] VDDI VSSI WL[1] S1AHSF400W40_MCB
XMCB_1<7> BL[7] BLB[7] VDDI VSSI WL[1] S1AHSF400W40_MCB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    ADR_X0_BIST_888
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ADR_X0_BIST_888 A[0] A[1] A[2] BIST1B BIST2 CK1B CK2 DEC_X0[0] 
+ DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] PD 
+ VDDHD VDDI VSSI XM[0] XM[1] XM[2]
*.PININFO A[0]:I A[1]:I A[2]:I BIST1B:I BIST2:I CK1B:I CK2:I PD:I XM[0]:I 
*.PININFO XM[1]:I XM[2]:I DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O 
*.PININFO DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O VDDHD:B VDDI:B VSSI:B
XI56<0> A[0] XM[0] AX[0] AXC[0] AXT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XI56<1> A[1] XM[1] AX[1] AXC[1] AXT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XI56<2> A[2] XM[2] AX[2] AXC[2] AXT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XIDEC_X0<0> NET11 NET11 DEC_X0[0] NET11 NET11 PD XA[0] VDDHD VSSI S1AHSF400W40_DECB1_X_SB
XIDEC_X0<1> NET11 NET11 DEC_X0[1] NET11 NET11 PD XA[1] VDDHD VSSI S1AHSF400W40_DECB1_X_SB
XIDEC_X0<2> NET11 NET11 DEC_X0[2] NET11 NET11 PD XA[2] VDDHD VSSI S1AHSF400W40_DECB1_X_SB
XIDEC_X0<3> NET11 NET11 DEC_X0[3] NET11 NET11 PD XA[3] VDDHD VSSI S1AHSF400W40_DECB1_X_SB
XIDEC_X0<4> NET11 NET11 DEC_X0[4] NET11 NET11 PD XA[4] VDDHD VSSI S1AHSF400W40_DECB1_X_SB
XIDEC_X0<5> NET11 NET11 DEC_X0[5] NET11 NET11 PD XA[5] VDDHD VSSI S1AHSF400W40_DECB1_X_SB
XIDEC_X0<6> NET11 NET11 DEC_X0[6] NET11 NET11 PD XA[6] VDDHD VSSI S1AHSF400W40_DECB1_X_SB
XIDEC_X0<7> NET11 NET11 DEC_X0[7] NET11 NET11 PD XA[7] VDDHD VSSI S1AHSF400W40_DECB1_X_SB
XI57<0> AXC[0] AXT[0] AXC[1] AXT[1] AXC[2] XA[0] XA[1] XA[2] XA[3] VDDHD VSSI 
+ S1AHSF400W40_DECB4_SB
XI57<1> AXC[0] AXT[0] AXC[1] AXT[1] AXT[2] XA[4] XA[5] XA[6] XA[7] VDDHD VSSI 
+ S1AHSF400W40_DECB4_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    ADR_X0_BIST_882
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ADR_X0_BIST_882 A[0] A[1] A[2] BIST1B BIST2 CK1B CK2 DEC_X0[0] 
+ DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] PD 
+ VDDHD VDDI VSSI XM[0] XM[1] XM[2]
*.PININFO A[0]:I A[1]:I A[2]:I BIST1B:I BIST2:I CK1B:I CK2:I PD:I XM[0]:I 
*.PININFO XM[1]:I XM[2]:I DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O 
*.PININFO DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O VDDHD:B VDDI:B VSSI:B
XI56<0> A[0] XM[0] AX[0] AXC[0] AXT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XI56<1> A[1] XM[1] AX[1] AXC[1] AXT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XI56<2> A[2] XM[2] AX[2] AXC[2] AXT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XIPDEC_X0<0> AXC[0] AXT[0] AXC[1] AXT[1] AXC[2] PD DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] VDDHD VSSI S1AHSF400W40_DECB4_882_SB
XIPDEC_X0<1> AXC[0] AXT[0] AXC[1] AXT[1] AXT[2] PD DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] VDDHD VSSI S1AHSF400W40_DECB4_882_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    ADR_X0_888
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ADR_X0_888 A[0] A[1] A[2] BIST1B BIST2 CK1B CK2 DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] PD VDDHD VDDI 
+ VSSI XM[0] XM[1] XM[2]
*.PININFO A[0]:I A[1]:I A[2]:I BIST1B:I BIST2:I CK1B:I CK2:I PD:I XM[0]:I 
*.PININFO XM[1]:I XM[2]:I DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O 
*.PININFO DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O VDDHD:B VDDI:B VSSI:B
XIDEC_X0<0> NET11 NET11 DEC_X0[0] NET11 NET11 PD XA[0] VDDHD VSSI S1AHSF400W40_DECB1_X_SB
XIDEC_X0<1> NET11 NET11 DEC_X0[1] NET11 NET11 PD XA[1] VDDHD VSSI S1AHSF400W40_DECB1_X_SB
XIDEC_X0<2> NET11 NET11 DEC_X0[2] NET11 NET11 PD XA[2] VDDHD VSSI S1AHSF400W40_DECB1_X_SB
XIDEC_X0<3> NET11 NET11 DEC_X0[3] NET11 NET11 PD XA[3] VDDHD VSSI S1AHSF400W40_DECB1_X_SB
XIDEC_X0<4> NET11 NET11 DEC_X0[4] NET11 NET11 PD XA[4] VDDHD VSSI S1AHSF400W40_DECB1_X_SB
XIDEC_X0<5> NET11 NET11 DEC_X0[5] NET11 NET11 PD XA[5] VDDHD VSSI S1AHSF400W40_DECB1_X_SB
XIDEC_X0<6> NET11 NET11 DEC_X0[6] NET11 NET11 PD XA[6] VDDHD VSSI S1AHSF400W40_DECB1_X_SB
XIDEC_X0<7> NET11 NET11 DEC_X0[7] NET11 NET11 PD XA[7] VDDHD VSSI S1AHSF400W40_DECB1_X_SB
XI57<0> AXC[0] AXT[0] AXC[1] AXT[1] AXC[2] XA[0] XA[1] XA[2] XA[3] VDDHD VSSI 
+ S1AHSF400W40_DECB4_SB
XI57<1> AXC[0] AXT[0] AXC[1] AXT[1] AXT[2] XA[4] XA[5] XA[6] XA[7] VDDHD VSSI 
+ S1AHSF400W40_DECB4_SB
XI56<0> A[0] XM[0] AX[0] AXC[0] AXT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XI56<1> A[1] XM[1] AX[1] AXC[1] AXT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XI56<2> A[2] XM[2] AX[2] AXC[2] AXT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    ADR_X0_882
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ADR_X0_882 A[0] A[1] A[2] BIST1B BIST2 CK1B CK2 DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] PD VDDHD VDDI 
+ VSSI XM[0] XM[1] XM[2]
*.PININFO A[0]:I A[1]:I A[2]:I BIST1B:I BIST2:I CK1B:I CK2:I PD:I XM[0]:I 
*.PININFO XM[1]:I XM[2]:I DEC_X0[0]:O DEC_X0[1]:O DEC_X0[2]:O DEC_X0[3]:O 
*.PININFO DEC_X0[4]:O DEC_X0[5]:O DEC_X0[6]:O DEC_X0[7]:O VDDHD:B VDDI:B VSSI:B
XI56<0> A[0] XM[0] AX[0] AXC[0] AXT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XI56<1> A[1] XM[1] AX[1] AXC[1] AXT[1] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XI56<2> A[2] XM[2] AX[2] AXC[2] AXT[2] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XIPDEC_X0<0> AXC[0] AXT[0] AXC[1] AXT[1] AXC[2] PD DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] VDDHD VSSI S1AHSF400W40_DECB4_882_SB
XIPDEC_X0<1> AXC[0] AXT[0] AXC[1] AXT[1] AXT[2] PD DEC_X0[4] DEC_X0[5] 
+ DEC_X0[6] DEC_X0[7] VDDHD VSSI S1AHSF400W40_DECB4_882_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    ADR_X2_BIST_888
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ADR_X2_BIST_888 A[0] A[1] A[2] BIST1B BIST2 CK1B CK2 CLK CLK_ENV 
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X2[4] DEC_X2[5] DEC_X2[6] 
+ DEC_X2[7] EN ENC PD VDDHD VDDI VSSI XM[0] XM[1] XM[2]
*.PININFO A[0]:I A[1]:I A[2]:I BIST1B:I BIST2:I CK1B:I CK2:I CLK:I CLK_ENV:I 
*.PININFO EN:I ENC:I PD:I XM[0]:I XM[1]:I XM[2]:I DEC_X2[0]:O DEC_X2[1]:O 
*.PININFO DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O DEC_X2[5]:O DEC_X2[6]:O 
*.PININFO DEC_X2[7]:O VDDHD:B VDDI:B VSSI:B
XI56<6> A[0] XM[0] AX[6] AXC[6] AXT[6] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XI56<7> A[1] XM[1] AX[7] AXC[7] AXT[7] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XI56<8> A[2] XM[2] AX[8] AXC[8] AXT[8] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XI54<0> AXC[6] AXT[6] AXC[7] AXT[7] AXC[8] XC[0] XC[1] XC[2] XC[3] VDDHD VSSI 
+ S1AHSF400W40_DECB4_SB
XI54<1> AXC[6] AXT[6] AXC[7] AXT[7] AXT[8] XC[4] XC[5] XC[6] XC[7] VDDHD VSSI 
+ S1AHSF400W40_DECB4_SB
XI55<0> CLK CLK_ENV DEC_X2[0] EN ENC PD XC[0] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XI55<1> CLK CLK_ENV DEC_X2[1] EN ENC PD XC[1] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XI55<2> CLK CLK_ENV DEC_X2[2] EN ENC PD XC[2] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XI55<3> CLK CLK_ENV DEC_X2[3] EN ENC PD XC[3] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XI55<4> CLK CLK_ENV DEC_X2[4] EN ENC PD XC[4] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XI55<5> CLK CLK_ENV DEC_X2[5] EN ENC PD XC[5] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XI55<6> CLK CLK_ENV DEC_X2[6] EN ENC PD XC[6] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XI55<7> CLK CLK_ENV DEC_X2[7] EN ENC PD XC[7] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    ADR_X2_BIST_884
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ADR_X2_BIST_884 A[0] A[1] BIST1B BIST2 CK1B CK2 CLK CLK_ENV DEC_X2[0] 
+ DEC_X2[1] DEC_X2[2] DEC_X2[3] EN ENC PD VDDHD VDDI VSSI XM[0] XM[1]
*.PININFO A[0]:I A[1]:I BIST1B:I BIST2:I CK1B:I CK2:I CLK:I CLK_ENV:I EN:I 
*.PININFO ENC:I PD:I XM[0]:I XM[1]:I DEC_X2[0]:O DEC_X2[1]:O DEC_X2[2]:O 
*.PININFO DEC_X2[3]:O VDDHD:B VDDI:B VSSI:B
XABUF_X<5> A[0] XM[0] AX[5] AXC[5] AXT[5] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XABUF_X<6> A[1] XM[1] AX[6] AXC[6] AXT[6] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XIDEC_X2<0> CLK CLK_ENV DEC_X2[0] EN ENC PD XC[0] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<1> CLK CLK_ENV DEC_X2[1] EN ENC PD XC[1] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<2> CLK CLK_ENV DEC_X2[2] EN ENC PD XC[2] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<3> CLK CLK_ENV DEC_X2[3] EN ENC PD XC[3] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIPDEC_X2<0> AXC[5] AXT[5] AXC[6] XC[0] XC[1] VDDHD VSSI S1AHSF400W40_DECB2_SB
XIPDEC_X2<1> AXC[5] AXT[5] AXT[6] XC[2] XC[3] VDDHD VSSI S1AHSF400W40_DECB2_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    ADR_X2_BIST_882
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ADR_X2_BIST_882 A[0] BIST1B BIST2 CK1B CK2 CLK CLK_ENV DEC_X2[0] 
+ DEC_X2[1] EN ENC PD VDDHD VDDI VSSI XM[0]
*.PININFO A[0]:I BIST1B:I BIST2:I CK1B:I CK2:I CLK:I CLK_ENV:I EN:I ENC:I PD:I 
*.PININFO XM[0]:I DEC_X2[0]:O DEC_X2[1]:O VDDHD:B VDDI:B VSSI:B
XABUF_X A[0] XM[0] AX[0] AXC[0] AXT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_BIST_SB
XIDEC_X2<0> CLK CLK_ENV DEC_X2[0] EN ENC PD AXC[0] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<1> CLK CLK_ENV DEC_X2[1] EN ENC PD AXT[0] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    ADR_X2_888
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ADR_X2_888 A[0] A[1] A[2] CK1B CK2 CLK CLK_ENV DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] DEC_X2[4] DEC_X2[5] DEC_X2[6] DEC_X2[7] EN ENC PD VDDHD 
+ VDDI VSSI
*.PININFO A[0]:I A[1]:I A[2]:I CK1B:I CK2:I CLK:I CLK_ENV:I EN:I ENC:I PD:I 
*.PININFO DEC_X2[0]:O DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O DEC_X2[4]:O 
*.PININFO DEC_X2[5]:O DEC_X2[6]:O DEC_X2[7]:O VDDHD:B VDDI:B VSSI:B
XI54<0> AXC[6] AXT[6] AXC[7] AXT[7] AXC[8] XC[0] XC[1] XC[2] XC[3] VDDHD VSSI 
+ S1AHSF400W40_DECB4_SB
XI54<1> AXC[6] AXT[6] AXC[7] AXT[7] AXT[8] XC[4] XC[5] XC[6] XC[7] VDDHD VSSI 
+ S1AHSF400W40_DECB4_SB
XI55<0> CLK CLK_ENV DEC_X2[0] EN ENC PD XC[0] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XI55<1> CLK CLK_ENV DEC_X2[1] EN ENC PD XC[1] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XI55<2> CLK CLK_ENV DEC_X2[2] EN ENC PD XC[2] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XI55<3> CLK CLK_ENV DEC_X2[3] EN ENC PD XC[3] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XI55<4> CLK CLK_ENV DEC_X2[4] EN ENC PD XC[4] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XI55<5> CLK CLK_ENV DEC_X2[5] EN ENC PD XC[5] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XI55<6> CLK CLK_ENV DEC_X2[6] EN ENC PD XC[6] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XI55<7> CLK CLK_ENV DEC_X2[7] EN ENC PD XC[7] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XI56<6> A[0] XM[6] AX[6] AXC[6] AXT[6] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XI56<7> A[1] XM[7] AX[7] AXC[7] AXT[7] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XI56<8> A[2] XM[8] AX[8] AXC[8] AXT[8] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    ADR_X2_884
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ADR_X2_884 A[0] A[1] CK1B CK2 CLK CLK_ENV DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] EN ENC PD VDDHD VDDI VSSI
*.PININFO A[0]:I A[1]:I CK1B:I CK2:I CLK:I CLK_ENV:I EN:I ENC:I PD:I 
*.PININFO DEC_X2[0]:O DEC_X2[1]:O DEC_X2[2]:O DEC_X2[3]:O VDDHD:B VDDI:B VSSI:B
XIDEC_X2<0> CLK CLK_ENV DEC_X2[0] EN ENC PD XC[0] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<1> CLK CLK_ENV DEC_X2[1] EN ENC PD XC[1] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<2> CLK CLK_ENV DEC_X2[2] EN ENC PD XC[2] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<3> CLK CLK_ENV DEC_X2[3] EN ENC PD XC[3] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XABUF_X<5> A[0] XM[5] AX[5] AXC[5] AXT[5] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XABUF_X<6> A[1] XM[6] AX[6] AXC[6] AXT[6] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_SB
XIPDEC_X2<0> AXC[5] AXT[5] AXC[6] XC[0] XC[1] VDDHD VSSI S1AHSF400W40_DECB2_SB
XIPDEC_X2<1> AXC[5] AXT[5] AXT[6] XC[2] XC[3] VDDHD VSSI S1AHSF400W40_DECB2_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    ADR_X2_882
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_ADR_X2_882 A[0] CK1B CK2 CLK CLK_ENV DEC_X2[0] DEC_X2[1] EN ENC PD 
+ VDDHD VDDI VSSI
*.PININFO A[0]:I CK1B:I CK2:I CLK:I CLK_ENV:I EN:I ENC:I PD:I DEC_X2[0]:O 
*.PININFO DEC_X2[1]:O VDDHD:B VDDI:B VSSI:B
XABUF_X A[0] XM[0] AX[0] AXC[0] AXT[0] BIST1B BIST2 CK1B CK2 VDDHD VSSI 
+ S1AHSF400W40_ABUF_882_SB
XIDEC_X2<0> CLK CLK_ENV DEC_X2[0] EN ENC PD AXC[0] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
XIDEC_X2<1> CLK CLK_ENV DEC_X2[1] EN ENC PD AXT[0] VDDHD VSSI S1AHSF400W40_DECB1_X2_SB
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MCNTIOX8_BIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCNTIOX8_BIST AWT BIST BLTRKWLDRV BWEB[0] BWEB[1] BWEB[2] BWEB[3] 
+ BWEB[4] BWEB[5] BWEB[6] BWEB[7] BWEBM[0] BWEBM[1] BWEBM[2] BWEBM[3] BWEBM[4] 
+ BWEBM[5] BWEBM[6] BWEBM[7] CEB CEBM CLK D[0] D[1] D[2] D[3] D[4] D[5] D[6] 
+ D[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] 
+ DM[0] DM[1] DM[2] DM[3] DM[4] DM[5] DM[6] DM[7] GBL[0] GBL[1] GBL[2] GBL[3] 
+ GBL[4] GBL[5] GBL[6] GBL[7] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] 
+ GBLB[6] GBLB[7] GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GWB[0] 
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] PD_BUF PD_CVDDBUF Q[0] Q[1] 
+ Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] REDEN REDENB RTSEL[0] RTSEL[1] RW_RE SLP TM 
+ TRKBL VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAE_TK WTSEL[0] WTSEL[1] 
+ WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] 
+ XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] 
+ YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I BWEB[0]:I BWEB[1]:I BWEB[2]:I BWEB[3]:I BWEB[4]:I 
*.PININFO BWEB[5]:I BWEB[6]:I BWEB[7]:I BWEBM[0]:I BWEBM[1]:I BWEBM[2]:I 
*.PININFO BWEBM[3]:I BWEBM[4]:I BWEBM[5]:I BWEBM[6]:I BWEBM[7]:I CEB:I CEBM:I 
*.PININFO CLK:I D[0]:I D[1]:I D[2]:I D[3]:I D[4]:I D[5]:I D[6]:I D[7]:I 
*.PININFO DM[0]:I DM[1]:I DM[2]:I DM[3]:I DM[4]:I DM[5]:I DM[6]:I DM[7]:I 
*.PININFO REDEN:I REDENB:I RTSEL[0]:I RTSEL[1]:I SLP:I TM:I WEB:I WEBM:I 
*.PININFO WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I 
*.PININFO X[5]:I X[6]:I X[7]:I X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I 
*.PININFO XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I 
*.PININFO Y[0]:I Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I Q[0]:O 
*.PININFO Q[1]:O Q[2]:O Q[3]:O Q[4]:O Q[5]:O Q[6]:O Q[7]:O VHI:O VLO:O 
*.PININFO BLTRKWLDRV:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B GBL[0]:B GBL[1]:B GBL[2]:B GBL[3]:B GBL[4]:B GBL[5]:B 
*.PININFO GBL[6]:B GBL[7]:B GBLB[0]:B GBLB[1]:B GBLB[2]:B GBLB[3]:B GBLB[4]:B 
*.PININFO GBLB[5]:B GBLB[6]:B GBLB[7]:B GW[0]:B GW[1]:B GW[2]:B GW[3]:B 
*.PININFO GW[4]:B GW[5]:B GW[6]:B GW[7]:B GWB[0]:B GWB[1]:B GWB[2]:B GWB[3]:B 
*.PININFO GWB[4]:B GWB[5]:B GWB[6]:B GWB[7]:B PD_BUF:B PD_CVDDBUF:B RW_RE:B 
*.PININFO TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XI8 AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] 
+ DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] SLP PD_BUF PD_CVDDBUF NET153 
+ REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL VDDHD VDDI VHI VLO VSSI WEB 
+ WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] 
+ X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] 
+ YM[3] S1AHSF400W40_CNT_CORE_M4_BIST
XIO_M8_L<0> AWT2 BIST2IO BWEB[0] BWEBM[0] CKD D[0] DM[0] GBL[0] GBLB[0] GW[0] 
+ GWB[0] PD_BUF Q[0] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XIO_M8_L<1> AWT2 BIST2IO BWEB[1] BWEBM[1] CKD D[1] DM[1] GBL[1] GBLB[1] GW[1] 
+ GWB[1] PD_BUF Q[1] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XIO_M8_L<2> AWT2 BIST2IO BWEB[2] BWEBM[2] CKD D[2] DM[2] GBL[2] GBLB[2] GW[2] 
+ GWB[2] PD_BUF Q[2] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XIO_M8_L<3> AWT2 BIST2IO BWEB[3] BWEBM[3] CKD D[3] DM[3] GBL[3] GBLB[3] GW[3] 
+ GWB[3] PD_BUF Q[3] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XI2<4> AWT2 BIST2IO BWEB[4] BWEBM[4] CKD D[4] DM[4] GBL[4] GBLB[4] GW[4] 
+ GWB[4] PD_BUF Q[4] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XI2<5> AWT2 BIST2IO BWEB[5] BWEBM[5] CKD D[5] DM[5] GBL[5] GBLB[5] GW[5] 
+ GWB[5] PD_BUF Q[5] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XI2<6> AWT2 BIST2IO BWEB[6] BWEBM[6] CKD D[6] DM[6] GBL[6] GBLB[6] GW[6] 
+ GWB[6] PD_BUF Q[6] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XI2<7> AWT2 BIST2IO BWEB[7] BWEBM[7] CKD D[7] DM[7] GBL[7] GBLB[7] GW[7] 
+ GWB[7] PD_BUF Q[7] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MCNTIOX2_BIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCNTIOX2_BIST AWT BIST BLTRKWLDRV BWEB[0] BWEB[1] BWEBM[0] BWEBM[1] 
+ CEB CEBM CLK D[0] D[1] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] 
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DM[0] DM[1] GBL[0] GBL[1] GBLB[0] GBLB[1] GW[0] GW[1] 
+ GWB[0] GWB[1] PD_BUF PD_CVDDBUF Q[0] Q[1] REDEN REDENB RTSEL[0] RTSEL[1] 
+ RW_RE SLP TM TRKBL VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] 
+ X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] 
+ Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I BWEB[0]:I BWEB[1]:I BWEBM[0]:I BWEBM[1]:I CEB:I CEBM:I 
*.PININFO CLK:I D[0]:I D[1]:I DM[0]:I DM[1]:I REDEN:I REDENB:I RTSEL[0]:I 
*.PININFO RTSEL[1]:I SLP:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I 
*.PININFO X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I 
*.PININFO X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I XM[5]:I 
*.PININFO XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I Y[2]:I Y[3]:I 
*.PININFO YM[0]:I YM[1]:I YM[2]:I YM[3]:I Q[0]:O Q[1]:O VHI:O VLO:O 
*.PININFO BLTRKWLDRV:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B GBL[0]:B GBL[1]:B GBLB[0]:B GBLB[1]:B GW[0]:B GW[1]:B 
*.PININFO GWB[0]:B GWB[1]:B PD_BUF:B PD_CVDDBUF:B RW_RE:B TRKBL:B VDDHD:B 
*.PININFO VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XI0 AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] 
+ DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] SLP PD_BUF PD_CVDDBUF NET86 
+ REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL VDDHD VDDI VHI VLO VSSI WEB 
+ WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] 
+ X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] 
+ YM[3] S1AHSF400W40_CNT_CORE_M16_BIST
XIO_M4_L AWT2 BIST2IO BWEB[0] BWEBM[0] CKD D[0] DM[0] GBL[0] GBLB[0] GW[0] 
+ GWB[0] PD_BUF Q[0] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M16
XI2 AWT2 BIST2IO BWEB[1] BWEBM[1] CKD D[1] DM[1] GBL[1] GBLB[1] GW[1] GWB[1] 
+ PD_BUF Q[1] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M16
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MCNTIOX4_BIST
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCNTIOX4_BIST AWT BIST BLTRKWLDRV BWEB[0] BWEB[1] BWEB[2] BWEB[3] 
+ BWEBM[0] BWEBM[1] BWEBM[2] BWEBM[3] CEB CEBM CLK D[0] D[1] D[2] D[3] 
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] 
+ DM[0] DM[1] DM[2] DM[3] GBL[0] GBL[1] GBL[2] GBL[3] GBLB[0] GBLB[1] GBLB[2] 
+ GBLB[3] GW[0] GW[1] GW[2] GW[3] GWB[0] GWB[1] GWB[2] GWB[3] PD_BUF 
+ PD_CVDDBUF Q[0] Q[1] Q[2] Q[3] REDEN REDENB RTSEL[0] RTSEL[1] RW_RE SLP TM 
+ TRKBL VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAE_TK WTSEL[0] WTSEL[1] 
+ WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] 
+ XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] 
+ YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I BWEB[0]:I BWEB[1]:I BWEB[2]:I BWEB[3]:I BWEBM[0]:I 
*.PININFO BWEBM[1]:I BWEBM[2]:I BWEBM[3]:I CEB:I CEBM:I CLK:I D[0]:I D[1]:I 
*.PININFO D[2]:I D[3]:I DM[0]:I DM[1]:I DM[2]:I DM[3]:I REDEN:I REDENB:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I SLP:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I 
*.PININFO XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I 
*.PININFO Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I Q[0]:O Q[1]:O Q[2]:O 
*.PININFO Q[3]:O VHI:O VLO:O BLTRKWLDRV:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B 
*.PININFO DEC_X0[3]:B DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B 
*.PININFO DEC_X1[0]:B DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B 
*.PININFO DEC_X1[5]:B DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B 
*.PININFO DEC_X2[2]:B DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B 
*.PININFO DEC_X3[3]:B DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B 
*.PININFO DEC_Y[0]:B DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B 
*.PININFO DEC_Y[6]:B DEC_Y[7]:B GBL[0]:B GBL[1]:B GBL[2]:B GBL[3]:B GBLB[0]:B 
*.PININFO GBLB[1]:B GBLB[2]:B GBLB[3]:B GW[0]:B GW[1]:B GW[2]:B GW[3]:B 
*.PININFO GWB[0]:B GWB[1]:B GWB[2]:B GWB[3]:B PD_BUF:B PD_CVDDBUF:B RW_RE:B 
*.PININFO TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XI7 AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] 
+ DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] SLP PD_BUF PD_CVDDBUF NET86 
+ REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL VDDHD VDDI VHI VLO VSSI WEB 
+ WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] 
+ X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] 
+ YM[3] S1AHSF400W40_CNT_CORE_M8_BIST
XIO_M8_L<0> AWT2 BIST2IO BWEB[0] BWEBM[0] CKD D[0] DM[0] GBL[0] GBLB[0] GW[0] 
+ GWB[0] PD_BUF Q[0] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M8
XIO_M8_L<1> AWT2 BIST2IO BWEB[1] BWEBM[1] CKD D[1] DM[1] GBL[1] GBLB[1] GW[1] 
+ GWB[1] PD_BUF Q[1] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M8
XI2<2> AWT2 BIST2IO BWEB[2] BWEBM[2] CKD D[2] DM[2] GBL[2] GBLB[2] GW[2] 
+ GWB[2] PD_BUF Q[2] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M8
XI2<3> AWT2 BIST2IO BWEB[3] BWEBM[3] CKD D[3] DM[3] GBL[3] GBLB[3] GW[3] 
+ GWB[3] PD_BUF Q[3] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M8
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LCTRL_F_M8_1S
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LCTRL_F_M8_1S BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] 
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] 
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] 
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF PD_CVDDBUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] 
+ WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE 
+ WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO DEC_Y[0]:I DEC_Y[1]:I DEC_Y[2]:I DEC_Y[3]:I DEC_Y[4]:I DEC_Y[5]:I 
*.PININFO DEC_Y[6]:I DEC_Y[7]:I PD_CVDDBUF:I YL[0]:I BLEQ_DN:O BLEQ_UP:O 
*.PININFO DEC_Y_DN[0]:O DEC_Y_DN[1]:O DEC_Y_DN[2]:O DEC_Y_DN[3]:O 
*.PININFO DEC_Y_DN[4]:O DEC_Y_DN[5]:O DEC_Y_DN[6]:O DEC_Y_DN[7]:O 
*.PININFO DEC_Y_UP[0]:O DEC_Y_UP[1]:O DEC_Y_UP[2]:O DEC_Y_UP[3]:O 
*.PININFO DEC_Y_UP[4]:O DEC_Y_UP[5]:O DEC_Y_UP[6]:O DEC_Y_UP[7]:O RE:O SAEB:O 
*.PININFO WE:O WLPY_DN[0]:O WLPY_DN[1]:O WLPY_DN[2]:O WLPY_DN[3]:O 
*.PININFO WLPY_UP[0]:O WLPY_UP[1]:O WLPY_UP[2]:O WLPY_UP[3]:O YL_LIO[0]:O 
*.PININFO YL_LIO[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B PD_BUF:B RW_RE:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B
XXDRV_WLP_D BLEQ_DN BLEQB_DN DEC_X3[0] PD_BUF WLP_SAE VDDHD VDDI VSSI 
+ WLPY_DN[0] S1AHSF400W40_XDRV_WLP_F
XLCNT BLEQB_DN BLEQB_UP DEC_X3[0] DEC_X3[1] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] 
+ DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] 
+ DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] 
+ DEC_Y_UP[6] DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLP_SAE 
+ YL[0] YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LCTRL_F_M16_1S
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LCTRL_F_M16_1S BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] 
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] 
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] 
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF PD_CVDDBUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] 
+ WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE 
+ WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO DEC_X2[0]:I DEC_X2[1]:I DEC_X2[2]:I DEC_X2[3]:I DEC_Y[0]:I 
*.PININFO DEC_Y[1]:I DEC_Y[2]:I DEC_Y[3]:I DEC_Y[4]:I DEC_Y[5]:I DEC_Y[6]:I 
*.PININFO DEC_Y[7]:I PD_BUF:I PD_CVDDBUF:I RW_RE:I WLP_SAE:I WLP_SAE_TK:I 
*.PININFO YL[0]:I BLEQ_DN:O BLEQ_UP:O DEC_Y_DN[0]:O DEC_Y_DN[1]:O 
*.PININFO DEC_Y_DN[2]:O DEC_Y_DN[3]:O DEC_Y_DN[4]:O DEC_Y_DN[5]:O 
*.PININFO DEC_Y_DN[6]:O DEC_Y_DN[7]:O DEC_Y_UP[0]:O DEC_Y_UP[1]:O 
*.PININFO DEC_Y_UP[2]:O DEC_Y_UP[3]:O DEC_Y_UP[4]:O DEC_Y_UP[5]:O 
*.PININFO DEC_Y_UP[6]:O DEC_Y_UP[7]:O RE:O SAEB:O WE:O WLPY_DN[0]:O 
*.PININFO WLPY_DN[1]:O WLPY_DN[2]:O WLPY_DN[3]:O WLPY_UP[0]:O WLPY_UP[1]:O 
*.PININFO WLPY_UP[2]:O WLPY_UP[3]:O YL_LIO[0]:O YL_LIO[1]:O DEC_X0[0]:B 
*.PININFO DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B DEC_X0[5]:B 
*.PININFO DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B DEC_X1[2]:B 
*.PININFO DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B DEC_X1[7]:B 
*.PININFO DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B DEC_X3[4]:B 
*.PININFO DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B VDDHD:B VDDI:B VSSI:B
XLCTRL_F_M8_1S BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] 
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] 
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] 
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF PD_CVDDBUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] 
+ WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE 
+ WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL_F_M8_1S
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LCTRL_F_M4_1S
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LCTRL_F_M4_1S BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] 
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] 
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] 
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF PD_CVDDBUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] 
+ WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE 
+ WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO DEC_Y[0]:I DEC_Y[1]:I DEC_Y[2]:I DEC_Y[3]:I DEC_Y[4]:I DEC_Y[5]:I 
*.PININFO DEC_Y[6]:I DEC_Y[7]:I PD_CVDDBUF:I YL[0]:I BLEQ_DN:O BLEQ_UP:O 
*.PININFO DEC_Y_DN[0]:O DEC_Y_DN[1]:O DEC_Y_DN[2]:O DEC_Y_DN[3]:O 
*.PININFO DEC_Y_DN[4]:O DEC_Y_DN[5]:O DEC_Y_DN[6]:O DEC_Y_DN[7]:O 
*.PININFO DEC_Y_UP[0]:O DEC_Y_UP[1]:O DEC_Y_UP[2]:O DEC_Y_UP[3]:O 
*.PININFO DEC_Y_UP[4]:O DEC_Y_UP[5]:O DEC_Y_UP[6]:O DEC_Y_UP[7]:O RE:O SAEB:O 
*.PININFO WE:O WLPY_DN[0]:O WLPY_DN[1]:O WLPY_DN[2]:O WLPY_DN[3]:O 
*.PININFO WLPY_UP[0]:O WLPY_UP[1]:O WLPY_UP[2]:O WLPY_UP[3]:O YL_LIO[0]:O 
*.PININFO YL_LIO[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B PD_BUF:B RW_RE:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B
XLCNT BLEQB_DN BLEQB_UP DEC_X3[0] DEC_X3[1] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] 
+ DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] 
+ DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] 
+ DEC_Y_UP[6] DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLP_SAE 
+ YL[0] YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL
XXDRV_WLP_D BLEQ_DN BLEQB_DN DEC_X3[0] PD_BUF WLP_SAE VDDHD VDDI VSSI 
+ WLPY_DN[0] S1AHSF400W40_XDRV_WLP_F
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LCTRL_S_M8_1S
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LCTRL_S_M8_1S BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] 
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] 
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] 
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF PD_CVDDBUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] 
+ WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE 
+ WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO DEC_Y[0]:I DEC_Y[1]:I DEC_Y[2]:I DEC_Y[3]:I DEC_Y[4]:I DEC_Y[5]:I 
*.PININFO DEC_Y[6]:I DEC_Y[7]:I PD_CVDDBUF:I YL[0]:I BLEQ_DN:O BLEQ_UP:O 
*.PININFO DEC_Y_DN[0]:O DEC_Y_DN[1]:O DEC_Y_DN[2]:O DEC_Y_DN[3]:O 
*.PININFO DEC_Y_DN[4]:O DEC_Y_DN[5]:O DEC_Y_DN[6]:O DEC_Y_DN[7]:O 
*.PININFO DEC_Y_UP[0]:O DEC_Y_UP[1]:O DEC_Y_UP[2]:O DEC_Y_UP[3]:O 
*.PININFO DEC_Y_UP[4]:O DEC_Y_UP[5]:O DEC_Y_UP[6]:O DEC_Y_UP[7]:O RE:O SAEB:O 
*.PININFO WE:O WLPY_DN[0]:O WLPY_DN[1]:O WLPY_DN[2]:O WLPY_DN[3]:O 
*.PININFO WLPY_UP[0]:O WLPY_UP[1]:O WLPY_UP[2]:O WLPY_UP[3]:O YL_LIO[0]:O 
*.PININFO YL_LIO[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B PD_BUF:B RW_RE:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B
XXDRV_WLP_DN BLEQ_DN BLEQB_DN DEC_X3[0] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] PD_BUF WLP_SAE VDDHD VDDI VSSI WLPY_DN[0] WLPY_DN[1] WLPY_DN[2] 
+ WLPY_DN[3] S1AHSF400W40_XDRV_WLP_S
XLCTRL BLEQB_DN BLEQB_UP DEC_X3[0] DEC_X3[1] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] 
+ DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] 
+ DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] 
+ DEC_Y_UP[6] DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLP_SAE 
+ YL[0] YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LCTRL_S_M16_1S
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LCTRL_S_M16_1S BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] 
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] 
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] 
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF PD_CVDDBUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] 
+ WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE 
+ WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO DEC_X2[0]:I DEC_X2[1]:I DEC_X2[2]:I DEC_X2[3]:I DEC_Y[0]:I 
*.PININFO DEC_Y[1]:I DEC_Y[2]:I DEC_Y[3]:I DEC_Y[4]:I DEC_Y[5]:I DEC_Y[6]:I 
*.PININFO DEC_Y[7]:I PD_BUF:I PD_CVDDBUF:I RW_RE:I WLP_SAE:I WLP_SAE_TK:I 
*.PININFO YL[0]:I BLEQ_DN:O BLEQ_UP:O DEC_Y_DN[0]:O DEC_Y_DN[1]:O 
*.PININFO DEC_Y_DN[2]:O DEC_Y_DN[3]:O DEC_Y_DN[4]:O DEC_Y_DN[5]:O 
*.PININFO DEC_Y_DN[6]:O DEC_Y_DN[7]:O DEC_Y_UP[0]:O DEC_Y_UP[1]:O 
*.PININFO DEC_Y_UP[2]:O DEC_Y_UP[3]:O DEC_Y_UP[4]:O DEC_Y_UP[5]:O 
*.PININFO DEC_Y_UP[6]:O DEC_Y_UP[7]:O RE:O SAEB:O WE:O WLPY_DN[0]:O 
*.PININFO WLPY_DN[1]:O WLPY_DN[2]:O WLPY_DN[3]:O WLPY_UP[0]:O WLPY_UP[1]:O 
*.PININFO WLPY_UP[2]:O WLPY_UP[3]:O YL_LIO[0]:O YL_LIO[1]:O DEC_X0[0]:B 
*.PININFO DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B DEC_X0[4]:B DEC_X0[5]:B 
*.PININFO DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B DEC_X1[1]:B DEC_X1[2]:B 
*.PININFO DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B DEC_X1[6]:B DEC_X1[7]:B 
*.PININFO DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B DEC_X3[4]:B 
*.PININFO DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B VDDHD:B VDDI:B VSSI:B
XLCTRL_S_M8_1S BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] 
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] 
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] 
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF PD_CVDDBUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] 
+ WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE 
+ WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL_S_M8_1S
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LCTRL_S_M4_1S
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LCTRL_S_M4_1S BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] 
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] 
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] 
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF PD_CVDDBUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] 
+ WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE 
+ WLP_SAE_TK YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO DEC_Y[0]:I DEC_Y[1]:I DEC_Y[2]:I DEC_Y[3]:I DEC_Y[4]:I DEC_Y[5]:I 
*.PININFO DEC_Y[6]:I DEC_Y[7]:I PD_CVDDBUF:I YL[0]:I BLEQ_DN:O BLEQ_UP:O 
*.PININFO DEC_Y_DN[0]:O DEC_Y_DN[1]:O DEC_Y_DN[2]:O DEC_Y_DN[3]:O 
*.PININFO DEC_Y_DN[4]:O DEC_Y_DN[5]:O DEC_Y_DN[6]:O DEC_Y_DN[7]:O 
*.PININFO DEC_Y_UP[0]:O DEC_Y_UP[1]:O DEC_Y_UP[2]:O DEC_Y_UP[3]:O 
*.PININFO DEC_Y_UP[4]:O DEC_Y_UP[5]:O DEC_Y_UP[6]:O DEC_Y_UP[7]:O RE:O SAEB:O 
*.PININFO WE:O WLPY_DN[0]:O WLPY_DN[1]:O WLPY_DN[2]:O WLPY_DN[3]:O 
*.PININFO WLPY_UP[0]:O WLPY_UP[1]:O WLPY_UP[2]:O WLPY_UP[3]:O YL_LIO[0]:O 
*.PININFO YL_LIO[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B PD_BUF:B RW_RE:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B
XLCTRL BLEQB_DN BLEQB_UP DEC_X3[0] DEC_X3[1] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] 
+ DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] 
+ DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] 
+ DEC_Y_UP[6] DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLP_SAE 
+ YL[0] YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL
XXDRV_WLP_DN BLEQ_DN BLEQB_DN DEC_X3[0] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] PD_BUF WLP_SAE VDDHD VDDI VSSI WLPY_DN[0] WLPY_DN[1] WLPY_DN[2] 
+ WLPY_DN[3] S1AHSF400W40_XDRV_WLP_S
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LIO_M16_1S
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LIO_M16_1S BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_DN[4] BLB_DN[5] 
+ BLB_DN[6] BLB_DN[7] BLB_DN[8] BLB_DN[9] BLB_DN[10] BLB_DN[11] BLB_DN[12] 
+ BLB_DN[13] BLB_DN[14] BLB_DN[15] BLB_UP[0] BLB_UP[1] BLB_UP[2] BLB_UP[3] 
+ BLB_UP[4] BLB_UP[5] BLB_UP[6] BLB_UP[7] BLB_UP[8] BLB_UP[9] BLB_UP[10] 
+ BLB_UP[11] BLB_UP[12] BLB_UP[13] BLB_UP[14] BLB_UP[15] BLEQ_DN BLEQ_UP 
+ BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] BL_DN[4] BL_DN[5] BL_DN[6] BL_DN[7] 
+ BL_DN[8] BL_DN[9] BL_DN[10] BL_DN[11] BL_DN[12] BL_DN[13] BL_DN[14] 
+ BL_DN[15] BL_UP[0] BL_UP[1] BL_UP[2] BL_UP[3] BL_UP[4] BL_UP[5] BL_UP[6] 
+ BL_UP[7] BL_UP[8] BL_UP[9] BL_UP[10] BL_UP[11] BL_UP[12] BL_UP[13] BL_UP[14] 
+ BL_UP[15] GBL GBLB GW GWB RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] 
+ Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] 
+ Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
*.PININFO BLEQ_DN:I BLEQ_UP:I GW:I GWB:I RE:I SAEB:I WE:I YL_LIO[0]:I 
*.PININFO YL_LIO[1]:I Y_DN[0]:I Y_DN[1]:I Y_DN[2]:I Y_DN[3]:I Y_DN[4]:I 
*.PININFO Y_DN[5]:I Y_DN[6]:I Y_DN[7]:I Y_UP[0]:I Y_UP[1]:I Y_UP[2]:I 
*.PININFO Y_UP[3]:I Y_UP[4]:I Y_UP[5]:I Y_UP[6]:I Y_UP[7]:I BLB_DN[0]:B 
*.PININFO BLB_DN[1]:B BLB_DN[2]:B BLB_DN[3]:B BLB_DN[4]:B BLB_DN[5]:B 
*.PININFO BLB_DN[6]:B BLB_DN[7]:B BLB_DN[8]:B BLB_DN[9]:B BLB_DN[10]:B 
*.PININFO BLB_DN[11]:B BLB_DN[12]:B BLB_DN[13]:B BLB_DN[14]:B BLB_DN[15]:B 
*.PININFO BLB_UP[0]:B BLB_UP[1]:B BLB_UP[2]:B BLB_UP[3]:B BLB_UP[4]:B 
*.PININFO BLB_UP[5]:B BLB_UP[6]:B BLB_UP[7]:B BLB_UP[8]:B BLB_UP[9]:B 
*.PININFO BLB_UP[10]:B BLB_UP[11]:B BLB_UP[12]:B BLB_UP[13]:B BLB_UP[14]:B 
*.PININFO BLB_UP[15]:B BL_DN[0]:B BL_DN[1]:B BL_DN[2]:B BL_DN[3]:B BL_DN[4]:B 
*.PININFO BL_DN[5]:B BL_DN[6]:B BL_DN[7]:B BL_DN[8]:B BL_DN[9]:B BL_DN[10]:B 
*.PININFO BL_DN[11]:B BL_DN[12]:B BL_DN[13]:B BL_DN[14]:B BL_DN[15]:B 
*.PININFO BL_UP[0]:B BL_UP[1]:B BL_UP[2]:B BL_UP[3]:B BL_UP[4]:B BL_UP[5]:B 
*.PININFO BL_UP[6]:B BL_UP[7]:B BL_UP[8]:B BL_UP[9]:B BL_UP[10]:B BL_UP[11]:B 
*.PININFO BL_UP[12]:B BL_UP[13]:B BL_UP[14]:B BL_UP[15]:B GBL:B GBLB:B VDDHD:B 
*.PININFO VDDI:B VSSI:B
XYPASS_DN_1 BL_DN[8] BL_DN[9] BL_DN[10] BL_DN[11] BL_DN[12] BL_DN[13] 
+ BL_DN[14] BL_DN[15] BLB_DN[8] BLB_DN[9] BLB_DN[10] BLB_DN[11] BLB_DN[12] 
+ BLB_DN[13] BLB_DN[14] BLB_DN[15] BLEQ_DN BLEQB_DN_1 DL_DN_1 DLB_DN_1 READ 
+ VDDI VSSI WC[1] WRITE WT[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] 
+ Y_DN[6] Y_DN[7] S1AHSF400W40_YPASS_M8
XYPASS_DN_0 BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] BL_DN[4] BL_DN[5] BL_DN[6] 
+ BL_DN[7] BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_DN[4] BLB_DN[5] 
+ BLB_DN[6] BLB_DN[7] BLEQ_DN BLEQB_DN_0 DL_DN_0 DLB_DN_0 READ VDDI VSSI WC[0] 
+ WRITE WT[0] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] 
+ S1AHSF400W40_YPASS_M8
XIO_RWBLK BLEQB_DN_0 BLEQB_DN_1 BLEQB_UP_0 BLEQB_UP_1 BLEQ_DN BLEQ_UP DLB_DN_0 
+ DLB_DN_1 DLB_UP_0 DLB_UP_1 DL_DN_0 DL_DN_1 DL_UP_0 DL_UP_1 GBL GBLB GW GWB 
+ RE READ SAEB VDDHD VDDI VSSI WC[0] WC[1] WE WRITE WT[0] WT[1] YL_LIO[0] 
+ YL_LIO[1] S1AHSF400W40_IO_RWBLK_M16
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LIO_M8_1S
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LIO_M8_1S BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_DN[4] BLB_DN[5] 
+ BLB_DN[6] BLB_DN[7] BLB_UP[0] BLB_UP[1] BLB_UP[2] BLB_UP[3] BLB_UP[4] 
+ BLB_UP[5] BLB_UP[6] BLB_UP[7] BLEQ_DN BLEQ_UP BL_DN[0] BL_DN[1] BL_DN[2] 
+ BL_DN[3] BL_DN[4] BL_DN[5] BL_DN[6] BL_DN[7] BL_UP[0] BL_UP[1] BL_UP[2] 
+ BL_UP[3] BL_UP[4] BL_UP[5] BL_UP[6] BL_UP[7] GBL GBLB GW GWB RE SAEB VDDHD 
+ VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] 
+ Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] 
+ Y_UP[6] Y_UP[7]
*.PININFO BLEQ_DN:I BLEQ_UP:I GW:I GWB:I RE:I SAEB:I WE:I YL_LIO[0]:I 
*.PININFO YL_LIO[1]:I Y_DN[0]:I Y_DN[1]:I Y_DN[2]:I Y_DN[3]:I Y_DN[4]:I 
*.PININFO Y_DN[5]:I Y_DN[6]:I Y_DN[7]:I Y_UP[0]:I Y_UP[1]:I Y_UP[2]:I 
*.PININFO Y_UP[3]:I Y_UP[4]:I Y_UP[5]:I Y_UP[6]:I Y_UP[7]:I BLB_DN[0]:B 
*.PININFO BLB_DN[1]:B BLB_DN[2]:B BLB_DN[3]:B BLB_DN[4]:B BLB_DN[5]:B 
*.PININFO BLB_DN[6]:B BLB_DN[7]:B BLB_UP[0]:B BLB_UP[1]:B BLB_UP[2]:B 
*.PININFO BLB_UP[3]:B BLB_UP[4]:B BLB_UP[5]:B BLB_UP[6]:B BLB_UP[7]:B 
*.PININFO BL_DN[0]:B BL_DN[1]:B BL_DN[2]:B BL_DN[3]:B BL_DN[4]:B BL_DN[5]:B 
*.PININFO BL_DN[6]:B BL_DN[7]:B BL_UP[0]:B BL_UP[1]:B BL_UP[2]:B BL_UP[3]:B 
*.PININFO BL_UP[4]:B BL_UP[5]:B BL_UP[6]:B BL_UP[7]:B GBL:B GBLB:B VDDHD:B 
*.PININFO VDDI:B VSSI:B
XIO_RWBLK BLEQB_DN_0 BLEQB_UP_0 BLEQ_DN BLEQ_UP DLB_DN DLB_UP DL_DN DL_UP GBL 
+ GBLB GW GWB RE READ SAEB VDDHD VDDI VSSI WC WE WRITE WT S1AHSF400W40_IO_RWBLK_M8
XYPASS_DN BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] BL_DN[4] BL_DN[5] BL_DN[6] 
+ BL_DN[7] BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_DN[4] BLB_DN[5] 
+ BLB_DN[6] BLB_DN[7] BLEQ_DN BLEQB_DN_0 DL_DN DLB_DN READ VDDI VSSI WC WRITE 
+ WT Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] S1AHSF400W40_YPASS_M8
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LIO_M4_1S
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LIO_M4_1S BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_UP[0] BLB_UP[1] 
+ BLB_UP[2] BLB_UP[3] BLEQ_DN BLEQ_UP BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] 
+ BL_UP[0] BL_UP[1] BL_UP[2] BL_UP[3] GBL GBLB GW GWB RE SAEB VDDHD VDDI VSSI 
+ WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] 
+ Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] 
+ Y_UP[7]
*.PININFO BLEQ_DN:I BLEQ_UP:I GW:I GWB:I RE:I SAEB:I WE:I YL_LIO[0]:I 
*.PININFO YL_LIO[1]:I Y_DN[0]:I Y_DN[1]:I Y_DN[2]:I Y_DN[3]:I Y_DN[4]:I 
*.PININFO Y_DN[5]:I Y_DN[6]:I Y_DN[7]:I Y_UP[0]:I Y_UP[1]:I Y_UP[2]:I 
*.PININFO Y_UP[3]:I Y_UP[4]:I Y_UP[5]:I Y_UP[6]:I Y_UP[7]:I BLB_DN[0]:B 
*.PININFO BLB_DN[1]:B BLB_DN[2]:B BLB_DN[3]:B BLB_UP[0]:B BLB_UP[1]:B 
*.PININFO BLB_UP[2]:B BLB_UP[3]:B BL_DN[0]:B BL_DN[1]:B BL_DN[2]:B BL_DN[3]:B 
*.PININFO BL_UP[0]:B BL_UP[1]:B BL_UP[2]:B BL_UP[3]:B GBL:B GBLB:B VDDHD:B 
*.PININFO VDDI:B VSSI:B
XIO_RWBLK BLEQB_DN_0 BLEQB_UP_0 BLEQ_DN BLEQ_UP DLB_DN DLB_UP DL_DN DL_UP GBL 
+ GBLB GW GWB SAEB VDDHD VDDI VSSI WC WT S1AHSF400W40_IO_RWBLK_M4
XYPASS_D BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] BLB_DN[0] BLB_DN[1] BLB_DN[2] 
+ BLB_DN[3] BLEQ_DN BLEQB_DN_0 DL_DN DLB_DN VDDI VSSI WC WT Y_DN[0] Y_DN[1] 
+ Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] S1AHSF400W40_YPASS_M4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MCNTIOX8
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCNTIOX8 AWT BIST BLTRKWLDRV BWEB[0] BWEB[1] BWEB[2] BWEB[3] BWEB[4] 
+ BWEB[5] BWEB[6] BWEB[7] BWEBM[0] BWEBM[1] BWEBM[2] BWEBM[3] BWEBM[4] 
+ BWEBM[5] BWEBM[6] BWEBM[7] CEB CEBM CLK D[0] D[1] D[2] D[3] D[4] D[5] D[6] 
+ D[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] 
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] 
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] 
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] 
+ DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] 
+ DM[0] DM[1] DM[2] DM[3] DM[4] DM[5] DM[6] DM[7] GBL[0] GBL[1] GBL[2] GBL[3] 
+ GBL[4] GBL[5] GBL[6] GBL[7] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] 
+ GBLB[6] GBLB[7] GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GWB[0] 
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] PD_BUF PD_CVDDBUF Q[0] Q[1] 
+ Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] REDEN REDENB RTSEL[0] RTSEL[1] RW_RE SLP TM 
+ TRKBL VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAE_TK WTSEL[0] WTSEL[1] 
+ WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] 
+ XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] 
+ YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I BWEB[0]:I BWEB[1]:I BWEB[2]:I BWEB[3]:I BWEB[4]:I 
*.PININFO BWEB[5]:I BWEB[6]:I BWEB[7]:I BWEBM[0]:I BWEBM[1]:I BWEBM[2]:I 
*.PININFO BWEBM[3]:I BWEBM[4]:I BWEBM[5]:I BWEBM[6]:I BWEBM[7]:I CEB:I CEBM:I 
*.PININFO CLK:I D[0]:I D[1]:I D[2]:I D[3]:I D[4]:I D[5]:I D[6]:I D[7]:I 
*.PININFO DM[0]:I DM[1]:I DM[2]:I DM[3]:I DM[4]:I DM[5]:I DM[6]:I DM[7]:I 
*.PININFO REDEN:I REDENB:I RTSEL[0]:I RTSEL[1]:I SLP:I TM:I WEB:I WEBM:I 
*.PININFO WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I 
*.PININFO X[5]:I X[6]:I X[7]:I X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I 
*.PININFO XM[3]:I XM[4]:I XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I 
*.PININFO Y[0]:I Y[1]:I Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I Q[0]:O 
*.PININFO Q[1]:O Q[2]:O Q[3]:O Q[4]:O Q[5]:O Q[6]:O Q[7]:O VHI:O VLO:O 
*.PININFO BLTRKWLDRV:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B GBL[0]:B GBL[1]:B GBL[2]:B GBL[3]:B GBL[4]:B GBL[5]:B 
*.PININFO GBL[6]:B GBL[7]:B GBLB[0]:B GBLB[1]:B GBLB[2]:B GBLB[3]:B GBLB[4]:B 
*.PININFO GBLB[5]:B GBLB[6]:B GBLB[7]:B GW[0]:B GW[1]:B GW[2]:B GW[3]:B 
*.PININFO GW[4]:B GW[5]:B GW[6]:B GW[7]:B GWB[0]:B GWB[1]:B GWB[2]:B GWB[3]:B 
*.PININFO GWB[4]:B GWB[5]:B GWB[6]:B GWB[7]:B PD_BUF:B PD_CVDDBUF:B RW_RE:B 
*.PININFO TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XI8 AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] 
+ DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] SLP PD_BUF PD_CVDDBUF NET153 
+ REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL VDDHD VDDI VHI VLO VSSI WEB 
+ WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] 
+ X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] 
+ YM[3] S1AHSF400W40_CNT_CORE_M4
XIO_M8_L<0> AWT2 BIST2IO BWEB[0] BWEBM[0] CKD D[0] DM[0] GBL[0] GBLB[0] GW[0] 
+ GWB[0] PD_BUF Q[0] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XIO_M8_L<1> AWT2 BIST2IO BWEB[1] BWEBM[1] CKD D[1] DM[1] GBL[1] GBLB[1] GW[1] 
+ GWB[1] PD_BUF Q[1] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XIO_M8_L<2> AWT2 BIST2IO BWEB[2] BWEBM[2] CKD D[2] DM[2] GBL[2] GBLB[2] GW[2] 
+ GWB[2] PD_BUF Q[2] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XIO_M8_L<3> AWT2 BIST2IO BWEB[3] BWEBM[3] CKD D[3] DM[3] GBL[3] GBLB[3] GW[3] 
+ GWB[3] PD_BUF Q[3] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XI2<4> AWT2 BIST2IO BWEB[4] BWEBM[4] CKD D[4] DM[4] GBL[4] GBLB[4] GW[4] 
+ GWB[4] PD_BUF Q[4] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XI2<5> AWT2 BIST2IO BWEB[5] BWEBM[5] CKD D[5] DM[5] GBL[5] GBLB[5] GW[5] 
+ GWB[5] PD_BUF Q[5] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XI2<6> AWT2 BIST2IO BWEB[6] BWEBM[6] CKD D[6] DM[6] GBL[6] GBLB[6] GW[6] 
+ GWB[6] PD_BUF Q[6] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
XI2<7> AWT2 BIST2IO BWEB[7] BWEBM[7] CKD D[7] DM[7] GBL[7] GBLB[7] GW[7] 
+ GWB[7] PD_BUF Q[7] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M4
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MCNTIOX4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCNTIOX4 AWT BIST BLTRKWLDRV BWEB[0] BWEB[1] BWEB[2] BWEB[3] BWEBM[0] 
+ BWEBM[1] BWEBM[2] BWEBM[3] CEB CEBM CLK D[0] D[1] D[2] D[3] DEC_X0[0] 
+ DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] 
+ DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] 
+ DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] 
+ DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] 
+ DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DM[0] DM[1] 
+ DM[2] DM[3] GBL[0] GBL[1] GBL[2] GBL[3] GBLB[0] GBLB[1] GBLB[2] GBLB[3] 
+ GW[0] GW[1] GW[2] GW[3] GWB[0] GWB[1] GWB[2] GWB[3] PD_BUF PD_CVDDBUF Q[0] 
+ Q[1] Q[2] Q[3] REDEN REDENB RTSEL[0] RTSEL[1] RW_RE SLP TM TRKBL VDDHD VDDI 
+ VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAE_TK WTSEL[0] WTSEL[1] WTSEL[2] X[0] 
+ X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] 
+ XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] 
+ YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I BWEB[0]:I BWEB[1]:I BWEB[2]:I BWEB[3]:I BWEBM[0]:I 
*.PININFO BWEBM[1]:I BWEBM[2]:I BWEBM[3]:I CEB:I CEBM:I CLK:I D[0]:I D[1]:I 
*.PININFO D[2]:I D[3]:I DM[0]:I DM[1]:I DM[2]:I DM[3]:I REDEN:I REDENB:I 
*.PININFO RTSEL[0]:I RTSEL[1]:I SLP:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I 
*.PININFO WTSEL[2]:I X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I 
*.PININFO X[8]:I X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I 
*.PININFO XM[5]:I XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I 
*.PININFO Y[2]:I Y[3]:I YM[0]:I YM[1]:I YM[2]:I YM[3]:I Q[0]:O Q[1]:O Q[2]:O 
*.PININFO Q[3]:O VHI:O VLO:O BLTRKWLDRV:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B 
*.PININFO DEC_X0[3]:B DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B 
*.PININFO DEC_X1[0]:B DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B 
*.PININFO DEC_X1[5]:B DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B 
*.PININFO DEC_X2[2]:B DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B 
*.PININFO DEC_X3[3]:B DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B 
*.PININFO DEC_Y[0]:B DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B 
*.PININFO DEC_Y[6]:B DEC_Y[7]:B GBL[0]:B GBL[1]:B GBL[2]:B GBL[3]:B GBLB[0]:B 
*.PININFO GBLB[1]:B GBLB[2]:B GBLB[3]:B GW[0]:B GW[1]:B GW[2]:B GW[3]:B 
*.PININFO GWB[0]:B GWB[1]:B GWB[2]:B GWB[3]:B PD_BUF:B PD_CVDDBUF:B RW_RE:B 
*.PININFO TRKBL:B VDDHD:B VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XI7 AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] 
+ DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] SLP PD_BUF PD_CVDDBUF NET86 
+ REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL VDDHD VDDI VHI VLO VSSI WEB 
+ WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] 
+ X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] 
+ YM[3] S1AHSF400W40_CNT_CORE_M8
XIO_M8_L<0> AWT2 BIST2IO BWEB[0] BWEBM[0] CKD D[0] DM[0] GBL[0] GBLB[0] GW[0] 
+ GWB[0] PD_BUF Q[0] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M8
XIO_M8_L<1> AWT2 BIST2IO BWEB[1] BWEBM[1] CKD D[1] DM[1] GBL[1] GBLB[1] GW[1] 
+ GWB[1] PD_BUF Q[1] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M8
XI2<2> AWT2 BIST2IO BWEB[2] BWEBM[2] CKD D[2] DM[2] GBL[2] GBLB[2] GW[2] 
+ GWB[2] PD_BUF Q[2] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M8
XI2<3> AWT2 BIST2IO BWEB[3] BWEBM[3] CKD D[3] DM[3] GBL[3] GBLB[3] GW[3] 
+ GWB[3] PD_BUF Q[3] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M8
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    TRKNOR
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TRKNOR BLB BLB_EDGE BL_EDGE BL_TK VDDI VSSI WL WL_TK TIEH
*.PININFO WL:I WL_TK:I TIEH:I BLB:B BLB_EDGE:B BL_EDGE:B BL_TK:B VDDI:B VSSI:B
XTKBL_EDGE BLB_EDGE BL_EDGE VDDI VSSI WL WL_TK TIEH S1AHSF400W40_TKBL_EDGE
XTKBL_BCELL BLB BL_TK VDDI VSSI WL WL_TK TIEH S1AHSF400W40_TKBL_BCELL
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    TRKNORX2
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TRKNORX2 BL_TK VDDI VSSI WL[0] WL[1] WL_TK FLOAT1 FLOAT2 FLOAT3 FLOAT4 
+ TIEH
*.PININFO WL[0]:I WL[1]:I WL_TK:I TIEH:I BL_TK:B VDDI:B VSSI:B FLOAT1:B 
*.PININFO FLOAT2:B FLOAT3:B FLOAT4:B
XTRKNOR_0 FLOAT4 FLOAT1 FLOAT3 BL_TK VDDI VSSI WL[0] WL_TK TIEH S1AHSF400W40_TRKNOR
XTRKNOR_1 FLOAT4 FLOAT1 FLOAT2 BL_TK VDDI VSSI WL[1] WL_TK TIEH S1AHSF400W40_TRKNOR
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MCB_TKWL_ISO
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCB_TKWL_ISO BL BLB VDDI VSSI WLL WLR
*.PININFO BL:B BLB:B VDDI:B VSSI:B WLL:B WLR:B
MNCHPD0 VSSI FLOAT_MCB BL_IN VSSI NCHPD_WISR L=0.065U W=0.140U M=1
MNCHPD1 BLB_IN FLOAT_MC VSSI VSSI NCHPD_WISR L=0.065U W=0.140U M=1
MPCHPU1 FLOAT_MCB FLOAT_MC VDDI VDDI PCHPU_WISR L=0.065U W=0.080U M=1
MPCHPU0 VDDI FLOAT_MCB FLOAT_MC VDDI PCHPU_WISR L=0.065U W=0.080U M=1
MNCHPG1 BLB WLR BLB_IN VSSI NCHPG_WISR L=0.075U W=0.090U M=1
MNCHPG0 BL_IN WLL BL VSSI NCHPG_WISR L=0.075U W=0.090U M=1
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    TKWL_2X2_ISO
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TKWL_2X2_ISO VDDI VSSI WL_TK_L[0] WL_TK_L[1] WL_TK_R[0] WL_TK_R[1]
*.PININFO WL_TK_L[0]:I WL_TK_L[1]:I WL_TK_R[0]:I WL_TK_R[1]:I VDDI:B VSSI:B
XTKWL_MCB_1 NET281 NET284 VDDI VSSI WL_TK_R[1] S1AHSF400W40_MCB_TKWL
XI24 NET030 NET284 VDDI VSSI WL_TK_R[0] S1AHSF400W40_MCB_TKWL
XI22 NET279 NET278 VDDI VSSI WL_TK_R[1] WL_TK_L[1] S1AHSF400W40_MCB_TKWL_ISO
XI25 NET294 NET278 VDDI VSSI WL_TK_R[0] WL_TK_L[0] S1AHSF400W40_MCB_TKWL_ISO
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    TKWL_ISO_X16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TKWL_ISO_X16 VDDI VSSI WL_TK_L[0] WL_TK_L[1] WL_TK_R[0] WL_TK_R[1]
*.PININFO VDDI:B VSSI:B WL_TK_L[0]:B WL_TK_L[1]:B WL_TK_R[0]:B WL_TK_R[1]:B
XI13 VDDI VSSI WL_TK_L[0] WL_TK_L[1] WL_TK_R[0] WL_TK_R[1] S1AHSF400W40_TKWL_2X2_ISO
XI14<0> VDDI VSSI WL_TK_R[0] WL_TK_R[1] S1AHSF400W40_TKWL_2X2
XI14<1> VDDI VSSI WL_TK_R[0] WL_TK_R[1] S1AHSF400W40_TKWL_2X2
XI14<2> VDDI VSSI WL_TK_R[0] WL_TK_R[1] S1AHSF400W40_TKWL_2X2
XI14<3> VDDI VSSI WL_TK_R[0] WL_TK_R[1] S1AHSF400W40_TKWL_2X2
XI14<4> VDDI VSSI WL_TK_R[0] WL_TK_R[1] S1AHSF400W40_TKWL_2X2
XI14<5> VDDI VSSI WL_TK_R[0] WL_TK_R[1] S1AHSF400W40_TKWL_2X2
XI14<6> VDDI VSSI WL_TK_R[0] WL_TK_R[1] S1AHSF400W40_TKWL_2X2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    TKWL_ISO_X8
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TKWL_ISO_X8 VDDI VSSI WL_TK_L[0] WL_TK_L[1] WL_TK_R[0] WL_TK_R[1]
*.PININFO VDDI:B VSSI:B WL_TK_L[0]:B WL_TK_L[1]:B WL_TK_R[0]:B WL_TK_R[1]:B
XI13 VDDI VSSI WL_TK_L[0] WL_TK_L[1] WL_TK_R[0] WL_TK_R[1] S1AHSF400W40_TKWL_2X2_ISO
XI14<0> VDDI VSSI WL_TK_R[0] WL_TK_R[1] S1AHSF400W40_TKWL_2X2
XI14<1> VDDI VSSI WL_TK_R[0] WL_TK_R[1] S1AHSF400W40_TKWL_2X2
XI14<2> VDDI VSSI WL_TK_R[0] WL_TK_R[1] S1AHSF400W40_TKWL_2X2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    TKWL_ISO_X4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TKWL_ISO_X4 VDDI VSSI WL_TK_L[0] WL_TK_L[1] WL_TK_R[0] WL_TK_R[1]
*.PININFO VDDI:B VSSI:B WL_TK_L[0]:B WL_TK_L[1]:B WL_TK_R[0]:B WL_TK_R[1]:B
XI13 VDDI VSSI WL_TK_L[0] WL_TK_L[1] WL_TK_R[0] WL_TK_R[1] S1AHSF400W40_TKWL_2X2_ISO
XI14 VDDI VSSI WL_TK_R[0] WL_TK_R[1] S1AHSF400W40_TKWL_2X2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    TKWL_2X16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TKWL_2X16 VDDI VSSI WL_DUM WL_TK
*.PININFO VDDI:B VSSI:B WL_DUM:B WL_TK:B
XI13<0> VDDI VSSI WL_DUM WL_TK S1AHSF400W40_TKWL_2X2
XI13<1> VDDI VSSI WL_DUM WL_TK S1AHSF400W40_TKWL_2X2
XI13<2> VDDI VSSI WL_DUM WL_TK S1AHSF400W40_TKWL_2X2
XI13<3> VDDI VSSI WL_DUM WL_TK S1AHSF400W40_TKWL_2X2
XI13<4> VDDI VSSI WL_DUM WL_TK S1AHSF400W40_TKWL_2X2
XI13<5> VDDI VSSI WL_DUM WL_TK S1AHSF400W40_TKWL_2X2
XI13<6> VDDI VSSI WL_DUM WL_TK S1AHSF400W40_TKWL_2X2
XI13<7> VDDI VSSI WL_DUM WL_TK S1AHSF400W40_TKWL_2X2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    TKWL_2X8
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TKWL_2X8 VDDI VSSI WL_DUM WL_TK
*.PININFO VDDI:B VSSI:B WL_DUM:B WL_TK:B
XI13<0> VDDI VSSI WL_DUM WL_TK S1AHSF400W40_TKWL_2X2
XI13<1> VDDI VSSI WL_DUM WL_TK S1AHSF400W40_TKWL_2X2
XI13<2> VDDI VSSI WL_DUM WL_TK S1AHSF400W40_TKWL_2X2
XI13<3> VDDI VSSI WL_DUM WL_TK S1AHSF400W40_TKWL_2X2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    TKWL_2X4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_TKWL_2X4 VDDI VSSI WL_DUM WL_TK
*.PININFO VDDI:B VSSI:B WL_DUM:B WL_TK:B
XI13 VDDI VSSI WL_DUM WL_TK S1AHSF400W40_TKWL_2X2
XI14 VDDI VSSI WL_DUM WL_TK S1AHSF400W40_TKWL_2X2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    MCNTIOX2
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_MCNTIOX2 AWT BIST BLTRKWLDRV BWEB[0] BWEB[1] BWEBM[0] BWEBM[1] CEB 
+ CEBM CLK D[0] D[1] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] 
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DM[0] DM[1] GBL[0] GBL[1] GBLB[0] GBLB[1] GW[0] GW[1] 
+ GWB[0] GWB[1] PD_BUF PD_CVDDBUF Q[0] Q[1] REDEN REDENB RTSEL[0] RTSEL[1] 
+ RW_RE SLP TM TRKBL VDDHD VDDI VHI VLO VSSI WEB WEBM WLP_SAE WLP_SAE_TK 
+ WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] X[3] X[4] X[5] X[6] X[7] X[8] X[9] 
+ X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] XM[6] XM[7] XM[8] XM[9] XM[10] 
+ Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] YM[3]
*.PININFO AWT:I BIST:I BWEB[0]:I BWEB[1]:I BWEBM[0]:I BWEBM[1]:I CEB:I CEBM:I 
*.PININFO CLK:I D[0]:I D[1]:I DM[0]:I DM[1]:I REDEN:I REDENB:I RTSEL[0]:I 
*.PININFO RTSEL[1]:I SLP:I TM:I WEB:I WEBM:I WTSEL[0]:I WTSEL[1]:I WTSEL[2]:I 
*.PININFO X[0]:I X[1]:I X[2]:I X[3]:I X[4]:I X[5]:I X[6]:I X[7]:I X[8]:I 
*.PININFO X[9]:I X[10]:I XM[0]:I XM[1]:I XM[2]:I XM[3]:I XM[4]:I XM[5]:I 
*.PININFO XM[6]:I XM[7]:I XM[8]:I XM[9]:I XM[10]:I Y[0]:I Y[1]:I Y[2]:I Y[3]:I 
*.PININFO YM[0]:I YM[1]:I YM[2]:I YM[3]:I Q[0]:O Q[1]:O VHI:O VLO:O 
*.PININFO BLTRKWLDRV:B DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B DEC_Y[0]:B 
*.PININFO DEC_Y[1]:B DEC_Y[2]:B DEC_Y[3]:B DEC_Y[4]:B DEC_Y[5]:B DEC_Y[6]:B 
*.PININFO DEC_Y[7]:B GBL[0]:B GBL[1]:B GBLB[0]:B GBLB[1]:B GW[0]:B GW[1]:B 
*.PININFO GWB[0]:B GWB[1]:B PD_BUF:B PD_CVDDBUF:B RW_RE:B TRKBL:B VDDHD:B 
*.PININFO VDDI:B VSSI:B WLP_SAE:B WLP_SAE_TK:B YL[0]:B
XIO_M4_L AWT2 BIST2IO BWEB[0] BWEBM[0] CKD D[0] DM[0] GBL[0] GBLB[0] GW[0] 
+ GWB[0] PD_BUF Q[0] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M16
XI2 AWT2 BIST2IO BWEB[1] BWEBM[1] CKD D[1] DM[1] GBL[1] GBLB[1] GW[1] GWB[1] 
+ PD_BUF Q[1] VDDHD VDDI VSSI WLP_SAEB S1AHSF400W40_IO_M16
XI0 AWT AWT2 BIST BIST2IO BLTRKWLDRV CEB CEBM CKD CLK DEC_X0[0] DEC_X0[1] 
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] 
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] 
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] 
+ DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] SLP PD_BUF PD_CVDDBUF NET86 
+ REDEN REDENB RTSEL[0] RTSEL[1] RW_RE TK TM TRKBL VDDHD VDDI VHI VLO VSSI WEB 
+ WEBM WLP_SAE WLP_SAEB WLP_SAE_TK WTSEL[0] WTSEL[1] WTSEL[2] X[0] X[1] X[2] 
+ X[3] X[4] X[5] X[6] X[7] X[8] X[9] X[10] XM[0] XM[1] XM[2] XM[3] XM[4] XM[5] 
+ XM[6] XM[7] XM[8] XM[9] XM[10] Y[0] Y[1] Y[2] Y[3] YL[0] YM[0] YM[1] YM[2] 
+ YM[3] S1AHSF400W40_CNT_CORE_M16
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    XDRV_WLP_M
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_XDRV_WLP_M BLEQ BLEQB BS DEC_X2[0] DEC_X2[1] PD_BUF RD_RST VDDHD VDDI 
+ VSSI WLOUT[0] WLOUT[1]
*.PININFO BS:I DEC_X2[0]:I DEC_X2[1]:I PD_BUF:I RD_RST:I BLEQ:O BLEQB:O 
*.PININFO WLOUT[0]:O WLOUT[1]:O VDDHD:B VDDI:B VSSI:B
MP6 SHARE RD_RSTB VDDHD VDDHD PCH L=60N W=780.0N M=1
MMP1115 NET268 NET212 VDDHD VDDHD PCH L=60N W=1.695U M=6
MP16 MWL2[0] DEC_X2[0] VDDHD VDDHD PCH L=60N W=360.0N M=1
MP20 BLEQB NET357 VDDHD VDDHD PCH L=60N W=2.25U M=4
MP18 MWL2[1] DEC_X2[1] VDDHD VDDHD PCH L=60N W=360.0N M=1
MP11 VDDHD RD_RSTB MWL2[1] VDDHD PCH L=60N W=750.0N M=2
MMP1114 WLOUT[0] NET244 VDDHD VDDHD PCH L=60N W=2.7U M=9
MP21 BLEQB BSB VDDHD VDDHD PCH L=60N W=2.25U M=4
MMP1112 WLOUT[1] NET268 VDDHD VDDHD PCH L=60N W=2.7U M=9
MP14 VDDHD RD_RSTB MWL2[0] VDDHD PCH L=60N W=750.0N M=2
MMP1118 NET244 NET216 VDDHD VDDHD PCH L=60N W=1.695U M=6
MN23 SHARE RD_RSTB VSSI VSSI NCH L=60N W=2.7U M=6
MMN1114 WLOUT[0] NET244 VSSI VSSI NCH L=60N W=2.265U M=6
MMN1118 NET244 NET216 VSSI VSSI NCH L=60N W=1.695U M=3
MN0 MWL2[0] DEC_X2[0] SHARE VSSI NCH L=60N W=750.0N M=2
MMN1115 NET268 NET212 VSSI VSSI NCH L=60N W=1.695U M=3
MMN1112 WLOUT[1] NET268 VSSI VSSI NCH L=60N W=2.265U M=6
MN18 BLEQB BSB NET264 VSSI NCH L=60N W=2.25U M=4
MN2 NET264 NET357 VSSI VSSI NCH L=60N W=2.25U M=4
MN6 MWL2[1] DEC_X2[1] SHARE VSSI NCH L=60N W=750.0N M=2
MN22 BLEQB PD_BUF VSSI VSSI NCH L=60N W=780.0N M=1
XNOR1 WLOUT[0] WLOUT[1] VSSI VDDHD NET357 S1AHSF400W40_ANOR FN2=1 WN2=0.2U LN2=0.1U FN1=1 
+ WN1=0.2U LN1=0.1U FP1=1 WP1=0.39U LP1=0.1U FP2=1 WP2=0.39U LP2=0.1U M=1
XI527 BSB RD_RST VSSI VDDHD RD_RSTB S1AHSF400W40_ANOR FN2=2 WN2=0.5U LN2=0.06U FN1=2 
+ WN1=0.5U LN1=0.06U FP1=2 WP1=1.5U LP1=0.06U FP2=2 WP2=1.5U LP2=0.06U M=1
XINV2 BLEQB VSSI VDDI BLEQ S1AHSF400W40_AINV FN=1 WN=1.5U LN=0.2U FP=1 WP=1.5U LP=0.2U 
+ M=18
XI497 MWL2[1] VSSI VDDHD NET212 S1AHSF400W40_AINV FN=1 WN=0.57U LN=0.2U FP=1 WP=1.125U 
+ LP=0.2U M=3
XINV21 MWL2[0] VSSI VDDHD NET216 S1AHSF400W40_AINV FN=1 WN=0.57U LN=0.2U FP=1 WP=1.125U 
+ LP=0.2U M=3
XI528 BS VSSI VDDHD BSB S1AHSF400W40_AINV FN=1 WN=0.5U LN=0.06U FP=1 WP=1U LP=0.06U M=2
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LCTRL_M_M8
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LCTRL_M_M8 BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] 
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] 
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] 
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF PD_CVDDBUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] 
+ WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE 
+ YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO DEC_Y[0]:I DEC_Y[1]:I DEC_Y[2]:I DEC_Y[3]:I DEC_Y[4]:I DEC_Y[5]:I 
*.PININFO DEC_Y[6]:I DEC_Y[7]:I PD_CVDDBUF:I YL[0]:I BLEQ_DN:O BLEQ_UP:O 
*.PININFO DEC_Y_DN[0]:O DEC_Y_DN[1]:O DEC_Y_DN[2]:O DEC_Y_DN[3]:O 
*.PININFO DEC_Y_DN[4]:O DEC_Y_DN[5]:O DEC_Y_DN[6]:O DEC_Y_DN[7]:O 
*.PININFO DEC_Y_UP[0]:O DEC_Y_UP[1]:O DEC_Y_UP[2]:O DEC_Y_UP[3]:O 
*.PININFO DEC_Y_UP[4]:O DEC_Y_UP[5]:O DEC_Y_UP[6]:O DEC_Y_UP[7]:O RE:O SAEB:O 
*.PININFO WE:O WLPY_DN[0]:O WLPY_DN[1]:O WLPY_DN[2]:O WLPY_DN[3]:O 
*.PININFO WLPY_UP[0]:O WLPY_UP[1]:O WLPY_UP[2]:O WLPY_UP[3]:O YL_LIO[0]:O 
*.PININFO YL_LIO[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B PD_BUF:B RW_RE:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE:B
XXDRV_WLP_UP BLEQ_UP BLEQB_UP DEC_X3[1] DEC_X2[0] DEC_X2[1] PD_BUF WLP_SAE 
+ VDDHD VDDI VSSI WLPY_UP[0] WLPY_UP[1] S1AHSF400W40_XDRV_WLP_M
XXDRV_WLP_DN BLEQ_DN BLEQB_DN DEC_X3[0] DEC_X2[0] DEC_X2[1] PD_BUF WLP_SAE 
+ VDDHD VDDI VSSI WLPY_DN[0] WLPY_DN[1] S1AHSF400W40_XDRV_WLP_M
XLCTRL BLEQB_DN BLEQB_UP DEC_X3[0] DEC_X3[1] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] 
+ DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] 
+ DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] 
+ DEC_Y_UP[6] DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLP_SAE 
+ YL[0] YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LCTRL_M_M16
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LCTRL_M_M16 BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] 
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] 
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] 
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF PD_CVDDBUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] 
+ WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE 
+ YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO DEC_X2[0]:I DEC_X2[1]:I DEC_X2[2]:I DEC_X2[3]:I DEC_Y[0]:I 
*.PININFO DEC_Y[1]:I DEC_Y[2]:I DEC_Y[3]:I DEC_Y[4]:I DEC_Y[5]:I DEC_Y[6]:I 
*.PININFO DEC_Y[7]:I PD_BUF:I PD_CVDDBUF:I RW_RE:I WLP_SAE:I YL[0]:I BLEQ_DN:O 
*.PININFO BLEQ_UP:O DEC_Y_DN[0]:O DEC_Y_DN[1]:O DEC_Y_DN[2]:O DEC_Y_DN[3]:O 
*.PININFO DEC_Y_DN[4]:O DEC_Y_DN[5]:O DEC_Y_DN[6]:O DEC_Y_DN[7]:O 
*.PININFO DEC_Y_UP[0]:O DEC_Y_UP[1]:O DEC_Y_UP[2]:O DEC_Y_UP[3]:O 
*.PININFO DEC_Y_UP[4]:O DEC_Y_UP[5]:O DEC_Y_UP[6]:O DEC_Y_UP[7]:O RE:O SAEB:O 
*.PININFO WE:O WLPY_DN[0]:O WLPY_DN[1]:O WLPY_DN[2]:O WLPY_DN[3]:O 
*.PININFO WLPY_UP[0]:O WLPY_UP[1]:O WLPY_UP[2]:O WLPY_UP[3]:O YL_LIO[0]:O 
*.PININFO YL_LIO[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B 
*.PININFO DEC_X3[3]:B DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B VDDHD:B 
*.PININFO VDDI:B VSSI:B
XLCTRL_M_M8 BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] 
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] 
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] 
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] 
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] 
+ DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF PD_CVDDBUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] 
+ WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE 
+ YL[0] YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL_M_M8
.ENDS

************************************************************************
* LIBRARY NAME: N65LP_SP_LEAFCELL
* CELL NAME:    LCTRL_M_M4
* VIEW NAME:    SCHEMATIC
************************************************************************

.SUBCKT S1AHSF400W40_LCTRL_M_M4 BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] 
+ DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] 
+ DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] 
+ DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] 
+ DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] 
+ DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] 
+ DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] 
+ DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] 
+ PD_BUF PD_CVDDBUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] 
+ WLPY_DN[2] WLPY_DN[3] WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE 
+ YL[0] YL_LIO[0] YL_LIO[1]
*.PININFO DEC_Y[0]:I DEC_Y[1]:I DEC_Y[2]:I DEC_Y[3]:I DEC_Y[4]:I DEC_Y[5]:I 
*.PININFO DEC_Y[6]:I DEC_Y[7]:I PD_CVDDBUF:I YL[0]:I BLEQ_DN:O BLEQ_UP:O 
*.PININFO DEC_Y_DN[0]:O DEC_Y_DN[1]:O DEC_Y_DN[2]:O DEC_Y_DN[3]:O 
*.PININFO DEC_Y_DN[4]:O DEC_Y_DN[5]:O DEC_Y_DN[6]:O DEC_Y_DN[7]:O 
*.PININFO DEC_Y_UP[0]:O DEC_Y_UP[1]:O DEC_Y_UP[2]:O DEC_Y_UP[3]:O 
*.PININFO DEC_Y_UP[4]:O DEC_Y_UP[5]:O DEC_Y_UP[6]:O DEC_Y_UP[7]:O RE:O SAEB:O 
*.PININFO WE:O WLPY_DN[0]:O WLPY_DN[1]:O WLPY_DN[2]:O WLPY_DN[3]:O 
*.PININFO WLPY_UP[0]:O WLPY_UP[1]:O WLPY_UP[2]:O WLPY_UP[3]:O YL_LIO[0]:O 
*.PININFO YL_LIO[1]:O DEC_X0[0]:B DEC_X0[1]:B DEC_X0[2]:B DEC_X0[3]:B 
*.PININFO DEC_X0[4]:B DEC_X0[5]:B DEC_X0[6]:B DEC_X0[7]:B DEC_X1[0]:B 
*.PININFO DEC_X1[1]:B DEC_X1[2]:B DEC_X1[3]:B DEC_X1[4]:B DEC_X1[5]:B 
*.PININFO DEC_X1[6]:B DEC_X1[7]:B DEC_X2[0]:B DEC_X2[1]:B DEC_X2[2]:B 
*.PININFO DEC_X2[3]:B DEC_X3[0]:B DEC_X3[1]:B DEC_X3[2]:B DEC_X3[3]:B 
*.PININFO DEC_X3[4]:B DEC_X3[5]:B DEC_X3[6]:B DEC_X3[7]:B PD_BUF:B RW_RE:B 
*.PININFO VDDHD:B VDDI:B VSSI:B WLP_SAE:B
XXDRV_WLP_UP BLEQ_UP BLEQB_UP DEC_X3[1] DEC_X2[0] DEC_X2[1] PD_BUF WLP_SAE 
+ VDDHD VDDI VSSI WLPY_UP[0] WLPY_UP[1] S1AHSF400W40_XDRV_WLP_M
XXDRV_WLP_DN BLEQ_DN BLEQB_DN DEC_X3[0] DEC_X2[0] DEC_X2[1] PD_BUF WLP_SAE 
+ VDDHD VDDI VSSI WLPY_DN[0] WLPY_DN[1] S1AHSF400W40_XDRV_WLP_M
XLCTRL BLEQB_DN BLEQB_UP DEC_X3[0] DEC_X3[1] DEC_Y[0] DEC_Y[1] DEC_Y[2] 
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] 
+ DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] 
+ DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] 
+ DEC_Y_UP[6] DEC_Y_UP[7] PD_BUF RE RW_RE SAEB VDDHD VDDI VSSI WE WLP_SAE 
+ YL[0] YL_LIO[0] YL_LIO[1] S1AHSF400W40_LCTRL
.ENDS




**** End of leaf cells

.SUBCKT S1AHSF400W40_CELL_ARR_X BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7]
+ BL[8] BL[9] BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18]
+ BL[19] BL[20] BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29]
+ BL[30] BL[31] BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40]
+ BL[41] BL[42] BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51]
+ BL[52] BL[53] BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62]
+ BL[63] BL[64] BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73]
+ BL[74] BL[75] BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84]
+ BL[85] BL[86] BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95]
+ BL[96] BL[97] BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105]
+ BL[106] BL[107] BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114]
+ BL[115] BL[116] BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123]
+ BL[124] BL[125] BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132]
+ BL[133] BL[134] BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141]
+ BL[142] BL[143] BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150]
+ BL[151] BL[152] BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159]
+ BL[160] BL[161] BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168]
+ BL[169] BL[170] BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177]
+ BL[178] BL[179] BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186]
+ BL[187] BL[188] BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195]
+ BL[196] BL[197] BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204]
+ BL[205] BL[206] BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213]
+ BL[214] BL[215] BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222]
+ BL[223] BL[224] BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231]
+ BL[232] BL[233] BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240]
+ BL[241] BL[242] BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249]
+ BL[250] BL[251] BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3]
+ BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13]
+ BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22]
+ BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31]
+ BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40]
+ BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49]
+ BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58]
+ BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67]
+ BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76]
+ BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85]
+ BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94]
+ BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103]
+ BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111]
+ BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119]
+ BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127]
+ BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135]
+ BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143]
+ BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151]
+ BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159]
+ BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167]
+ BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175]
+ BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183]
+ BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191]
+ BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199]
+ BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207]
+ BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215]
+ BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223]
+ BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231]
+ BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239]
+ BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247]
+ BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[0]
+ WL[1] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8]
+ GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18]
+ GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27]
+ GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36]
+ GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45]
+ GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54]
+ GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63]
+ GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8]
+ GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16]
+ GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24]
+ GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32]
+ GBLB[33] GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40]
+ GBLB[41] GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48]
+ GBLB[49] GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56]
+ GBLB[57] GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1]
+ GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13]
+ GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24]
+ GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35]
+ GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46]
+ GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57]
+ GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4]
+ GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14]
+ GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23]
+ GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32]
+ GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41]
+ GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50]
+ GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59]
+ GWB[60] GWB[61] GWB[62] GWB[63]
XMCB_0 BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] GBL[0] GBLB[0] GW[0]
+ GWB[0] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_1 BL[4] BL[5] BL[6] BL[7] BLB[4] BLB[5] BLB[6] BLB[7] GBL[1] GBLB[1] GW[1]
+ GWB[1] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_2 BL[8] BL[9] BL[10] BL[11] BLB[8] BLB[9] BLB[10] BLB[11] GBL[2] GBLB[2]
+ GW[2] GWB[2] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_3 BL[12] BL[13] BL[14] BL[15] BLB[12] BLB[13] BLB[14] BLB[15] GBL[3]
+ GBLB[3] GW[3] GWB[3] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_4 BL[16] BL[17] BL[18] BL[19] BLB[16] BLB[17] BLB[18] BLB[19] GBL[4]
+ GBLB[4] GW[4] GWB[4] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_5 BL[20] BL[21] BL[22] BL[23] BLB[20] BLB[21] BLB[22] BLB[23] GBL[5]
+ GBLB[5] GW[5] GWB[5] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_6 BL[24] BL[25] BL[26] BL[27] BLB[24] BLB[25] BLB[26] BLB[27] GBL[6]
+ GBLB[6] GW[6] GWB[6] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_7 BL[28] BL[29] BL[30] BL[31] BLB[28] BLB[29] BLB[30] BLB[31] GBL[7]
+ GBLB[7] GW[7] GWB[7] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_8 BL[32] BL[33] BL[34] BL[35] BLB[32] BLB[33] BLB[34] BLB[35] GBL[8]
+ GBLB[8] GW[8] GWB[8] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_9 BL[36] BL[37] BL[38] BL[39] BLB[36] BLB[37] BLB[38] BLB[39] GBL[9]
+ GBLB[9] GW[9] GWB[9] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_10 BL[40] BL[41] BL[42] BL[43] BLB[40] BLB[41] BLB[42] BLB[43] GBL[10]
+ GBLB[10] GW[10] GWB[10] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_11 BL[44] BL[45] BL[46] BL[47] BLB[44] BLB[45] BLB[46] BLB[47] GBL[11]
+ GBLB[11] GW[11] GWB[11] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_12 BL[48] BL[49] BL[50] BL[51] BLB[48] BLB[49] BLB[50] BLB[51] GBL[12]
+ GBLB[12] GW[12] GWB[12] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_13 BL[52] BL[53] BL[54] BL[55] BLB[52] BLB[53] BLB[54] BLB[55] GBL[13]
+ GBLB[13] GW[13] GWB[13] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_14 BL[56] BL[57] BL[58] BL[59] BLB[56] BLB[57] BLB[58] BLB[59] GBL[14]
+ GBLB[14] GW[14] GWB[14] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_15 BL[60] BL[61] BL[62] BL[63] BLB[60] BLB[61] BLB[62] BLB[63] GBL[15]
+ GBLB[15] GW[15] GWB[15] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_16 BL[64] BL[65] BL[66] BL[67] BLB[64] BLB[65] BLB[66] BLB[67] GBL[16]
+ GBLB[16] GW[16] GWB[16] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_17 BL[68] BL[69] BL[70] BL[71] BLB[68] BLB[69] BLB[70] BLB[71] GBL[17]
+ GBLB[17] GW[17] GWB[17] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_18 BL[72] BL[73] BL[74] BL[75] BLB[72] BLB[73] BLB[74] BLB[75] GBL[18]
+ GBLB[18] GW[18] GWB[18] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_19 BL[76] BL[77] BL[78] BL[79] BLB[76] BLB[77] BLB[78] BLB[79] GBL[19]
+ GBLB[19] GW[19] GWB[19] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_20 BL[80] BL[81] BL[82] BL[83] BLB[80] BLB[81] BLB[82] BLB[83] GBL[20]
+ GBLB[20] GW[20] GWB[20] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_21 BL[84] BL[85] BL[86] BL[87] BLB[84] BLB[85] BLB[86] BLB[87] GBL[21]
+ GBLB[21] GW[21] GWB[21] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_22 BL[88] BL[89] BL[90] BL[91] BLB[88] BLB[89] BLB[90] BLB[91] GBL[22]
+ GBLB[22] GW[22] GWB[22] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_23 BL[92] BL[93] BL[94] BL[95] BLB[92] BLB[93] BLB[94] BLB[95] GBL[23]
+ GBLB[23] GW[23] GWB[23] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_24 BL[96] BL[97] BL[98] BL[99] BLB[96] BLB[97] BLB[98] BLB[99] GBL[24]
+ GBLB[24] GW[24] GWB[24] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_25 BL[100] BL[101] BL[102] BL[103] BLB[100] BLB[101] BLB[102] BLB[103]
+ GBL[25] GBLB[25] GW[25] GWB[25] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_26 BL[104] BL[105] BL[106] BL[107] BLB[104] BLB[105] BLB[106] BLB[107]
+ GBL[26] GBLB[26] GW[26] GWB[26] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_27 BL[108] BL[109] BL[110] BL[111] BLB[108] BLB[109] BLB[110] BLB[111]
+ GBL[27] GBLB[27] GW[27] GWB[27] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_28 BL[112] BL[113] BL[114] BL[115] BLB[112] BLB[113] BLB[114] BLB[115]
+ GBL[28] GBLB[28] GW[28] GWB[28] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_29 BL[116] BL[117] BL[118] BL[119] BLB[116] BLB[117] BLB[118] BLB[119]
+ GBL[29] GBLB[29] GW[29] GWB[29] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_30 BL[120] BL[121] BL[122] BL[123] BLB[120] BLB[121] BLB[122] BLB[123]
+ GBL[30] GBLB[30] GW[30] GWB[30] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_31 BL[124] BL[125] BL[126] BL[127] BLB[124] BLB[125] BLB[126] BLB[127]
+ GBL[31] GBLB[31] GW[31] GWB[31] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_32 BL[128] BL[129] BL[130] BL[131] BLB[128] BLB[129] BLB[130] BLB[131]
+ GBL[32] GBLB[32] GW[32] GWB[32] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_33 BL[132] BL[133] BL[134] BL[135] BLB[132] BLB[133] BLB[134] BLB[135]
+ GBL[33] GBLB[33] GW[33] GWB[33] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_34 BL[136] BL[137] BL[138] BL[139] BLB[136] BLB[137] BLB[138] BLB[139]
+ GBL[34] GBLB[34] GW[34] GWB[34] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_35 BL[140] BL[141] BL[142] BL[143] BLB[140] BLB[141] BLB[142] BLB[143]
+ GBL[35] GBLB[35] GW[35] GWB[35] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_36 BL[144] BL[145] BL[146] BL[147] BLB[144] BLB[145] BLB[146] BLB[147]
+ GBL[36] GBLB[36] GW[36] GWB[36] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_37 BL[148] BL[149] BL[150] BL[151] BLB[148] BLB[149] BLB[150] BLB[151]
+ GBL[37] GBLB[37] GW[37] GWB[37] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_38 BL[152] BL[153] BL[154] BL[155] BLB[152] BLB[153] BLB[154] BLB[155]
+ GBL[38] GBLB[38] GW[38] GWB[38] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_39 BL[156] BL[157] BL[158] BL[159] BLB[156] BLB[157] BLB[158] BLB[159]
+ GBL[39] GBLB[39] GW[39] GWB[39] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_40 BL[160] BL[161] BL[162] BL[163] BLB[160] BLB[161] BLB[162] BLB[163]
+ GBL[40] GBLB[40] GW[40] GWB[40] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_41 BL[164] BL[165] BL[166] BL[167] BLB[164] BLB[165] BLB[166] BLB[167]
+ GBL[41] GBLB[41] GW[41] GWB[41] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_42 BL[168] BL[169] BL[170] BL[171] BLB[168] BLB[169] BLB[170] BLB[171]
+ GBL[42] GBLB[42] GW[42] GWB[42] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_43 BL[172] BL[173] BL[174] BL[175] BLB[172] BLB[173] BLB[174] BLB[175]
+ GBL[43] GBLB[43] GW[43] GWB[43] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_44 BL[176] BL[177] BL[178] BL[179] BLB[176] BLB[177] BLB[178] BLB[179]
+ GBL[44] GBLB[44] GW[44] GWB[44] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_45 BL[180] BL[181] BL[182] BL[183] BLB[180] BLB[181] BLB[182] BLB[183]
+ GBL[45] GBLB[45] GW[45] GWB[45] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_46 BL[184] BL[185] BL[186] BL[187] BLB[184] BLB[185] BLB[186] BLB[187]
+ GBL[46] GBLB[46] GW[46] GWB[46] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_47 BL[188] BL[189] BL[190] BL[191] BLB[188] BLB[189] BLB[190] BLB[191]
+ GBL[47] GBLB[47] GW[47] GWB[47] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_48 BL[192] BL[193] BL[194] BL[195] BLB[192] BLB[193] BLB[194] BLB[195]
+ GBL[48] GBLB[48] GW[48] GWB[48] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_49 BL[196] BL[197] BL[198] BL[199] BLB[196] BLB[197] BLB[198] BLB[199]
+ GBL[49] GBLB[49] GW[49] GWB[49] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_50 BL[200] BL[201] BL[202] BL[203] BLB[200] BLB[201] BLB[202] BLB[203]
+ GBL[50] GBLB[50] GW[50] GWB[50] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_51 BL[204] BL[205] BL[206] BL[207] BLB[204] BLB[205] BLB[206] BLB[207]
+ GBL[51] GBLB[51] GW[51] GWB[51] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_52 BL[208] BL[209] BL[210] BL[211] BLB[208] BLB[209] BLB[210] BLB[211]
+ GBL[52] GBLB[52] GW[52] GWB[52] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_53 BL[212] BL[213] BL[214] BL[215] BLB[212] BLB[213] BLB[214] BLB[215]
+ GBL[53] GBLB[53] GW[53] GWB[53] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_54 BL[216] BL[217] BL[218] BL[219] BLB[216] BLB[217] BLB[218] BLB[219]
+ GBL[54] GBLB[54] GW[54] GWB[54] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_55 BL[220] BL[221] BL[222] BL[223] BLB[220] BLB[221] BLB[222] BLB[223]
+ GBL[55] GBLB[55] GW[55] GWB[55] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_56 BL[224] BL[225] BL[226] BL[227] BLB[224] BLB[225] BLB[226] BLB[227]
+ GBL[56] GBLB[56] GW[56] GWB[56] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_57 BL[228] BL[229] BL[230] BL[231] BLB[228] BLB[229] BLB[230] BLB[231]
+ GBL[57] GBLB[57] GW[57] GWB[57] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_58 BL[232] BL[233] BL[234] BL[235] BLB[232] BLB[233] BLB[234] BLB[235]
+ GBL[58] GBLB[58] GW[58] GWB[58] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_59 BL[236] BL[237] BL[238] BL[239] BLB[236] BLB[237] BLB[238] BLB[239]
+ GBL[59] GBLB[59] GW[59] GWB[59] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_60 BL[240] BL[241] BL[242] BL[243] BLB[240] BLB[241] BLB[242] BLB[243]
+ GBL[60] GBLB[60] GW[60] GWB[60] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_61 BL[244] BL[245] BL[246] BL[247] BLB[244] BLB[245] BLB[246] BLB[247]
+ GBL[61] GBLB[61] GW[61] GWB[61] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_62 BL[248] BL[249] BL[250] BL[251] BLB[248] BLB[249] BLB[250] BLB[251]
+ GBL[62] GBLB[62] GW[62] GWB[62] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
XMCB_63 BL[252] BL[253] BL[254] BL[255] BLB[252] BLB[253] BLB[254] BLB[255]
+ GBL[63] GBLB[63] GW[63] GWB[63] VDDI VSSI WL[0] WL[1] S1AHSF400W40_MCB_2X4
.ENDS

.SUBCKT S1AHSF400W40_CELL_ARR_XY_F BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6]
+ BL[7] BL[8] BL[9] BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17]
+ BL[18] BL[19] BL[20] BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28]
+ BL[29] BL[30] BL[31] BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39]
+ BL[40] BL[41] BL[42] BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50]
+ BL[51] BL[52] BL[53] BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61]
+ BL[62] BL[63] BL[64] BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72]
+ BL[73] BL[74] BL[75] BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83]
+ BL[84] BL[85] BL[86] BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94]
+ BL[95] BL[96] BL[97] BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104]
+ BL[105] BL[106] BL[107] BL[108] BL[109] BL[110] BL[111] BL[112] BL[113]
+ BL[114] BL[115] BL[116] BL[117] BL[118] BL[119] BL[120] BL[121] BL[122]
+ BL[123] BL[124] BL[125] BL[126] BL[127] BL[128] BL[129] BL[130] BL[131]
+ BL[132] BL[133] BL[134] BL[135] BL[136] BL[137] BL[138] BL[139] BL[140]
+ BL[141] BL[142] BL[143] BL[144] BL[145] BL[146] BL[147] BL[148] BL[149]
+ BL[150] BL[151] BL[152] BL[153] BL[154] BL[155] BL[156] BL[157] BL[158]
+ BL[159] BL[160] BL[161] BL[162] BL[163] BL[164] BL[165] BL[166] BL[167]
+ BL[168] BL[169] BL[170] BL[171] BL[172] BL[173] BL[174] BL[175] BL[176]
+ BL[177] BL[178] BL[179] BL[180] BL[181] BL[182] BL[183] BL[184] BL[185]
+ BL[186] BL[187] BL[188] BL[189] BL[190] BL[191] BL[192] BL[193] BL[194]
+ BL[195] BL[196] BL[197] BL[198] BL[199] BL[200] BL[201] BL[202] BL[203]
+ BL[204] BL[205] BL[206] BL[207] BL[208] BL[209] BL[210] BL[211] BL[212]
+ BL[213] BL[214] BL[215] BL[216] BL[217] BL[218] BL[219] BL[220] BL[221]
+ BL[222] BL[223] BL[224] BL[225] BL[226] BL[227] BL[228] BL[229] BL[230]
+ BL[231] BL[232] BL[233] BL[234] BL[235] BL[236] BL[237] BL[238] BL[239]
+ BL[240] BL[241] BL[242] BL[243] BL[244] BL[245] BL[246] BL[247] BL[248]
+ BL[249] BL[250] BL[251] BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2]
+ BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12]
+ BLB[13] BLB[14] BLB[15] BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21]
+ BLB[22] BLB[23] BLB[24] BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30]
+ BLB[31] BLB[32] BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39]
+ BLB[40] BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48]
+ BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57]
+ BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66]
+ BLB[67] BLB[68] BLB[69] BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75]
+ BLB[76] BLB[77] BLB[78] BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84]
+ BLB[85] BLB[86] BLB[87] BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93]
+ BLB[94] BLB[95] BLB[96] BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102]
+ BLB[103] BLB[104] BLB[105] BLB[106] BLB[107] BLB[108] BLB[109] BLB[110]
+ BLB[111] BLB[112] BLB[113] BLB[114] BLB[115] BLB[116] BLB[117] BLB[118]
+ BLB[119] BLB[120] BLB[121] BLB[122] BLB[123] BLB[124] BLB[125] BLB[126]
+ BLB[127] BLB[128] BLB[129] BLB[130] BLB[131] BLB[132] BLB[133] BLB[134]
+ BLB[135] BLB[136] BLB[137] BLB[138] BLB[139] BLB[140] BLB[141] BLB[142]
+ BLB[143] BLB[144] BLB[145] BLB[146] BLB[147] BLB[148] BLB[149] BLB[150]
+ BLB[151] BLB[152] BLB[153] BLB[154] BLB[155] BLB[156] BLB[157] BLB[158]
+ BLB[159] BLB[160] BLB[161] BLB[162] BLB[163] BLB[164] BLB[165] BLB[166]
+ BLB[167] BLB[168] BLB[169] BLB[170] BLB[171] BLB[172] BLB[173] BLB[174]
+ BLB[175] BLB[176] BLB[177] BLB[178] BLB[179] BLB[180] BLB[181] BLB[182]
+ BLB[183] BLB[184] BLB[185] BLB[186] BLB[187] BLB[188] BLB[189] BLB[190]
+ BLB[191] BLB[192] BLB[193] BLB[194] BLB[195] BLB[196] BLB[197] BLB[198]
+ BLB[199] BLB[200] BLB[201] BLB[202] BLB[203] BLB[204] BLB[205] BLB[206]
+ BLB[207] BLB[208] BLB[209] BLB[210] BLB[211] BLB[212] BLB[213] BLB[214]
+ BLB[215] BLB[216] BLB[217] BLB[218] BLB[219] BLB[220] BLB[221] BLB[222]
+ BLB[223] BLB[224] BLB[225] BLB[226] BLB[227] BLB[228] BLB[229] BLB[230]
+ BLB[231] BLB[232] BLB[233] BLB[234] BLB[235] BLB[236] BLB[237] BLB[238]
+ BLB[239] BLB[240] BLB[241] BLB[242] BLB[243] BLB[244] BLB[245] BLB[246]
+ BLB[247] BLB[248] BLB[249] BLB[250] BLB[251] BLB[252] BLB[253] BLB[254]
+ BLB[255] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10]
+ WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21]
+ WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32]
+ WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43]
+ WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54]
+ WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63]
XCELL_ARR_X_0 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6]
+ BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15] BLB[16]
+ BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24] BLB[25]
+ BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33] BLB[34]
+ BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42] BLB[43]
+ BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51] BLB[52]
+ BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60] BLB[61]
+ BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69] BLB[70]
+ BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78] BLB[79]
+ BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87] BLB[88]
+ BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96] BLB[97]
+ BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105] BLB[106]
+ BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113] BLB[114]
+ BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121] BLB[122]
+ BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129] BLB[130]
+ BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137] BLB[138]
+ BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145] BLB[146]
+ BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153] BLB[154]
+ BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161] BLB[162]
+ BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169] BLB[170]
+ BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177] BLB[178]
+ BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185] BLB[186]
+ BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193] BLB[194]
+ BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201] BLB[202]
+ BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209] BLB[210]
+ BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217] BLB[218]
+ BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225] BLB[226]
+ BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233] BLB[234]
+ BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241] BLB[242]
+ BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249] BLB[250]
+ BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[0] WL[1] VDDI VSSI GBL[0]
+ GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11]
+ GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20]
+ GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29]
+ GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38]
+ GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47]
+ GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56]
+ GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3] GW[4]
+ GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16]
+ GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27]
+ GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37] GW[38]
+ GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48] GW[49]
+ GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59] GW[60]
+ GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7]
+ GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17]
+ GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26]
+ GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35]
+ GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44]
+ GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53]
+ GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62]
+ GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_1 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6]
+ BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15] BLB[16]
+ BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24] BLB[25]
+ BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33] BLB[34]
+ BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42] BLB[43]
+ BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51] BLB[52]
+ BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60] BLB[61]
+ BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69] BLB[70]
+ BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78] BLB[79]
+ BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87] BLB[88]
+ BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96] BLB[97]
+ BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105] BLB[106]
+ BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113] BLB[114]
+ BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121] BLB[122]
+ BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129] BLB[130]
+ BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137] BLB[138]
+ BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145] BLB[146]
+ BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153] BLB[154]
+ BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161] BLB[162]
+ BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169] BLB[170]
+ BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177] BLB[178]
+ BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185] BLB[186]
+ BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193] BLB[194]
+ BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201] BLB[202]
+ BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209] BLB[210]
+ BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217] BLB[218]
+ BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225] BLB[226]
+ BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233] BLB[234]
+ BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241] BLB[242]
+ BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249] BLB[250]
+ BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[2] WL[3] VDDI VSSI GBL[0]
+ GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11]
+ GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20]
+ GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29]
+ GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38]
+ GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47]
+ GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56]
+ GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3] GW[4]
+ GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16]
+ GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27]
+ GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37] GW[38]
+ GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48] GW[49]
+ GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59] GW[60]
+ GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7]
+ GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17]
+ GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26]
+ GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35]
+ GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44]
+ GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53]
+ GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62]
+ GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_2 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6]
+ BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15] BLB[16]
+ BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24] BLB[25]
+ BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33] BLB[34]
+ BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42] BLB[43]
+ BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51] BLB[52]
+ BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60] BLB[61]
+ BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69] BLB[70]
+ BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78] BLB[79]
+ BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87] BLB[88]
+ BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96] BLB[97]
+ BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105] BLB[106]
+ BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113] BLB[114]
+ BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121] BLB[122]
+ BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129] BLB[130]
+ BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137] BLB[138]
+ BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145] BLB[146]
+ BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153] BLB[154]
+ BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161] BLB[162]
+ BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169] BLB[170]
+ BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177] BLB[178]
+ BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185] BLB[186]
+ BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193] BLB[194]
+ BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201] BLB[202]
+ BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209] BLB[210]
+ BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217] BLB[218]
+ BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225] BLB[226]
+ BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233] BLB[234]
+ BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241] BLB[242]
+ BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249] BLB[250]
+ BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[4] WL[5] VDDI VSSI GBL[0]
+ GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11]
+ GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20]
+ GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29]
+ GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38]
+ GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47]
+ GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56]
+ GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3] GW[4]
+ GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16]
+ GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27]
+ GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37] GW[38]
+ GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48] GW[49]
+ GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59] GW[60]
+ GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7]
+ GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17]
+ GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26]
+ GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35]
+ GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44]
+ GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53]
+ GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62]
+ GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_3 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6]
+ BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15] BLB[16]
+ BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24] BLB[25]
+ BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33] BLB[34]
+ BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42] BLB[43]
+ BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51] BLB[52]
+ BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60] BLB[61]
+ BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69] BLB[70]
+ BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78] BLB[79]
+ BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87] BLB[88]
+ BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96] BLB[97]
+ BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105] BLB[106]
+ BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113] BLB[114]
+ BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121] BLB[122]
+ BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129] BLB[130]
+ BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137] BLB[138]
+ BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145] BLB[146]
+ BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153] BLB[154]
+ BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161] BLB[162]
+ BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169] BLB[170]
+ BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177] BLB[178]
+ BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185] BLB[186]
+ BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193] BLB[194]
+ BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201] BLB[202]
+ BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209] BLB[210]
+ BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217] BLB[218]
+ BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225] BLB[226]
+ BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233] BLB[234]
+ BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241] BLB[242]
+ BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249] BLB[250]
+ BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[6] WL[7] VDDI VSSI GBL[0]
+ GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11]
+ GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20]
+ GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29]
+ GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38]
+ GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47]
+ GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56]
+ GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3] GW[4]
+ GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16]
+ GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27]
+ GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37] GW[38]
+ GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48] GW[49]
+ GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59] GW[60]
+ GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7]
+ GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17]
+ GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26]
+ GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35]
+ GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44]
+ GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53]
+ GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62]
+ GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_4 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6]
+ BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15] BLB[16]
+ BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24] BLB[25]
+ BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33] BLB[34]
+ BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42] BLB[43]
+ BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51] BLB[52]
+ BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60] BLB[61]
+ BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69] BLB[70]
+ BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78] BLB[79]
+ BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87] BLB[88]
+ BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96] BLB[97]
+ BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105] BLB[106]
+ BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113] BLB[114]
+ BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121] BLB[122]
+ BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129] BLB[130]
+ BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137] BLB[138]
+ BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145] BLB[146]
+ BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153] BLB[154]
+ BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161] BLB[162]
+ BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169] BLB[170]
+ BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177] BLB[178]
+ BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185] BLB[186]
+ BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193] BLB[194]
+ BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201] BLB[202]
+ BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209] BLB[210]
+ BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217] BLB[218]
+ BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225] BLB[226]
+ BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233] BLB[234]
+ BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241] BLB[242]
+ BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249] BLB[250]
+ BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[8] WL[9] VDDI VSSI GBL[0]
+ GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11]
+ GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20]
+ GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29]
+ GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38]
+ GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47]
+ GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56]
+ GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3] GW[4]
+ GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16]
+ GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27]
+ GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37] GW[38]
+ GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48] GW[49]
+ GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59] GW[60]
+ GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7]
+ GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17]
+ GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26]
+ GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35]
+ GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44]
+ GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53]
+ GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62]
+ GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_5 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6]
+ BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15] BLB[16]
+ BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24] BLB[25]
+ BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33] BLB[34]
+ BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42] BLB[43]
+ BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51] BLB[52]
+ BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60] BLB[61]
+ BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69] BLB[70]
+ BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78] BLB[79]
+ BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87] BLB[88]
+ BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96] BLB[97]
+ BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105] BLB[106]
+ BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113] BLB[114]
+ BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121] BLB[122]
+ BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129] BLB[130]
+ BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137] BLB[138]
+ BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145] BLB[146]
+ BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153] BLB[154]
+ BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161] BLB[162]
+ BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169] BLB[170]
+ BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177] BLB[178]
+ BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185] BLB[186]
+ BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193] BLB[194]
+ BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201] BLB[202]
+ BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209] BLB[210]
+ BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217] BLB[218]
+ BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225] BLB[226]
+ BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233] BLB[234]
+ BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241] BLB[242]
+ BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249] BLB[250]
+ BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[10] WL[11] VDDI VSSI GBL[0]
+ GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11]
+ GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20]
+ GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29]
+ GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38]
+ GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47]
+ GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56]
+ GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3] GW[4]
+ GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16]
+ GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27]
+ GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37] GW[38]
+ GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48] GW[49]
+ GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59] GW[60]
+ GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7]
+ GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17]
+ GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26]
+ GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35]
+ GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44]
+ GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53]
+ GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62]
+ GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_6 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6]
+ BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15] BLB[16]
+ BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24] BLB[25]
+ BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33] BLB[34]
+ BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42] BLB[43]
+ BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51] BLB[52]
+ BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60] BLB[61]
+ BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69] BLB[70]
+ BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78] BLB[79]
+ BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87] BLB[88]
+ BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96] BLB[97]
+ BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105] BLB[106]
+ BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113] BLB[114]
+ BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121] BLB[122]
+ BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129] BLB[130]
+ BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137] BLB[138]
+ BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145] BLB[146]
+ BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153] BLB[154]
+ BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161] BLB[162]
+ BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169] BLB[170]
+ BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177] BLB[178]
+ BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185] BLB[186]
+ BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193] BLB[194]
+ BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201] BLB[202]
+ BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209] BLB[210]
+ BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217] BLB[218]
+ BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225] BLB[226]
+ BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233] BLB[234]
+ BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241] BLB[242]
+ BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249] BLB[250]
+ BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[12] WL[13] VDDI VSSI GBL[0]
+ GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11]
+ GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20]
+ GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29]
+ GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38]
+ GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47]
+ GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56]
+ GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3] GW[4]
+ GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16]
+ GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27]
+ GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37] GW[38]
+ GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48] GW[49]
+ GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59] GW[60]
+ GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7]
+ GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17]
+ GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26]
+ GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35]
+ GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44]
+ GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53]
+ GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62]
+ GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_7 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6]
+ BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15] BLB[16]
+ BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24] BLB[25]
+ BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33] BLB[34]
+ BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42] BLB[43]
+ BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51] BLB[52]
+ BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60] BLB[61]
+ BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69] BLB[70]
+ BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78] BLB[79]
+ BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87] BLB[88]
+ BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96] BLB[97]
+ BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105] BLB[106]
+ BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113] BLB[114]
+ BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121] BLB[122]
+ BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129] BLB[130]
+ BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137] BLB[138]
+ BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145] BLB[146]
+ BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153] BLB[154]
+ BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161] BLB[162]
+ BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169] BLB[170]
+ BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177] BLB[178]
+ BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185] BLB[186]
+ BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193] BLB[194]
+ BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201] BLB[202]
+ BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209] BLB[210]
+ BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217] BLB[218]
+ BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225] BLB[226]
+ BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233] BLB[234]
+ BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241] BLB[242]
+ BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249] BLB[250]
+ BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[14] WL[15] VDDI VSSI GBL[0]
+ GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11]
+ GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20]
+ GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29]
+ GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38]
+ GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47]
+ GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56]
+ GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3] GW[4]
+ GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16]
+ GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27]
+ GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37] GW[38]
+ GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48] GW[49]
+ GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59] GW[60]
+ GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7]
+ GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17]
+ GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26]
+ GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35]
+ GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44]
+ GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53]
+ GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62]
+ GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_8 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6]
+ BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15] BLB[16]
+ BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24] BLB[25]
+ BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33] BLB[34]
+ BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42] BLB[43]
+ BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51] BLB[52]
+ BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60] BLB[61]
+ BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69] BLB[70]
+ BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78] BLB[79]
+ BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87] BLB[88]
+ BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96] BLB[97]
+ BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105] BLB[106]
+ BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113] BLB[114]
+ BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121] BLB[122]
+ BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129] BLB[130]
+ BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137] BLB[138]
+ BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145] BLB[146]
+ BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153] BLB[154]
+ BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161] BLB[162]
+ BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169] BLB[170]
+ BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177] BLB[178]
+ BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185] BLB[186]
+ BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193] BLB[194]
+ BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201] BLB[202]
+ BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209] BLB[210]
+ BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217] BLB[218]
+ BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225] BLB[226]
+ BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233] BLB[234]
+ BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241] BLB[242]
+ BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249] BLB[250]
+ BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[16] WL[17] VDDI VSSI GBL[0]
+ GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11]
+ GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20]
+ GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29]
+ GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38]
+ GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47]
+ GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56]
+ GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3] GW[4]
+ GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16]
+ GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27]
+ GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37] GW[38]
+ GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48] GW[49]
+ GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59] GW[60]
+ GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7]
+ GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17]
+ GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26]
+ GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35]
+ GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44]
+ GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53]
+ GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62]
+ GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_9 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9] BL[10]
+ BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21]
+ BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BL[32]
+ BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42] BL[43]
+ BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54]
+ BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64] BL[65]
+ BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75] BL[76]
+ BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86] BL[87]
+ BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97] BL[98]
+ BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107] BL[108]
+ BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116] BL[117]
+ BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125] BL[126]
+ BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134] BL[135]
+ BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143] BL[144]
+ BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152] BL[153]
+ BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161] BL[162]
+ BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170] BL[171]
+ BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179] BL[180]
+ BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188] BL[189]
+ BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197] BL[198]
+ BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206] BL[207]
+ BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215] BL[216]
+ BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224] BL[225]
+ BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233] BL[234]
+ BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242] BL[243]
+ BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251] BL[252]
+ BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5] BLB[6]
+ BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15] BLB[16]
+ BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24] BLB[25]
+ BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33] BLB[34]
+ BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42] BLB[43]
+ BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51] BLB[52]
+ BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60] BLB[61]
+ BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69] BLB[70]
+ BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78] BLB[79]
+ BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87] BLB[88]
+ BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96] BLB[97]
+ BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105] BLB[106]
+ BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113] BLB[114]
+ BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121] BLB[122]
+ BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129] BLB[130]
+ BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137] BLB[138]
+ BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145] BLB[146]
+ BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153] BLB[154]
+ BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161] BLB[162]
+ BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169] BLB[170]
+ BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177] BLB[178]
+ BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185] BLB[186]
+ BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193] BLB[194]
+ BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201] BLB[202]
+ BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209] BLB[210]
+ BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217] BLB[218]
+ BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225] BLB[226]
+ BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233] BLB[234]
+ BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241] BLB[242]
+ BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249] BLB[250]
+ BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[18] WL[19] VDDI VSSI GBL[0]
+ GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11]
+ GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19] GBL[20]
+ GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28] GBL[29]
+ GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37] GBL[38]
+ GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46] GBL[47]
+ GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55] GBL[56]
+ GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0] GBLB[1]
+ GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10]
+ GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17] GBLB[18]
+ GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25] GBLB[26]
+ GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33] GBLB[34]
+ GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41] GBLB[42]
+ GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49] GBLB[50]
+ GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57] GBLB[58]
+ GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3] GW[4]
+ GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16]
+ GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27]
+ GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37] GW[38]
+ GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48] GW[49]
+ GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59] GW[60]
+ GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7]
+ GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17]
+ GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26]
+ GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35]
+ GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44]
+ GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53]
+ GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62]
+ GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_10 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[20] WL[21] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_11 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[22] WL[23] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_12 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[24] WL[25] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_13 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[26] WL[27] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_14 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[28] WL[29] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_15 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[30] WL[31] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_16 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[32] WL[33] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_17 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[34] WL[35] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_18 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[36] WL[37] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_19 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[38] WL[39] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_20 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[40] WL[41] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_21 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[42] WL[43] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_22 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[44] WL[45] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_23 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[46] WL[47] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_24 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[48] WL[49] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_25 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[50] WL[51] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_26 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[52] WL[53] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_27 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[54] WL[55] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_28 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[56] WL[57] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_29 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[58] WL[59] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_30 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[60] WL[61] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
XCELL_ARR_X_31 BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8] BL[9]
+ BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BL[16] BL[17] BL[18] BL[19] BL[20]
+ BL[21] BL[22] BL[23] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31]
+ BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BL[40] BL[41] BL[42]
+ BL[43] BL[44] BL[45] BL[46] BL[47] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53]
+ BL[54] BL[55] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BL[64]
+ BL[65] BL[66] BL[67] BL[68] BL[69] BL[70] BL[71] BL[72] BL[73] BL[74] BL[75]
+ BL[76] BL[77] BL[78] BL[79] BL[80] BL[81] BL[82] BL[83] BL[84] BL[85] BL[86]
+ BL[87] BL[88] BL[89] BL[90] BL[91] BL[92] BL[93] BL[94] BL[95] BL[96] BL[97]
+ BL[98] BL[99] BL[100] BL[101] BL[102] BL[103] BL[104] BL[105] BL[106] BL[107]
+ BL[108] BL[109] BL[110] BL[111] BL[112] BL[113] BL[114] BL[115] BL[116]
+ BL[117] BL[118] BL[119] BL[120] BL[121] BL[122] BL[123] BL[124] BL[125]
+ BL[126] BL[127] BL[128] BL[129] BL[130] BL[131] BL[132] BL[133] BL[134]
+ BL[135] BL[136] BL[137] BL[138] BL[139] BL[140] BL[141] BL[142] BL[143]
+ BL[144] BL[145] BL[146] BL[147] BL[148] BL[149] BL[150] BL[151] BL[152]
+ BL[153] BL[154] BL[155] BL[156] BL[157] BL[158] BL[159] BL[160] BL[161]
+ BL[162] BL[163] BL[164] BL[165] BL[166] BL[167] BL[168] BL[169] BL[170]
+ BL[171] BL[172] BL[173] BL[174] BL[175] BL[176] BL[177] BL[178] BL[179]
+ BL[180] BL[181] BL[182] BL[183] BL[184] BL[185] BL[186] BL[187] BL[188]
+ BL[189] BL[190] BL[191] BL[192] BL[193] BL[194] BL[195] BL[196] BL[197]
+ BL[198] BL[199] BL[200] BL[201] BL[202] BL[203] BL[204] BL[205] BL[206]
+ BL[207] BL[208] BL[209] BL[210] BL[211] BL[212] BL[213] BL[214] BL[215]
+ BL[216] BL[217] BL[218] BL[219] BL[220] BL[221] BL[222] BL[223] BL[224]
+ BL[225] BL[226] BL[227] BL[228] BL[229] BL[230] BL[231] BL[232] BL[233]
+ BL[234] BL[235] BL[236] BL[237] BL[238] BL[239] BL[240] BL[241] BL[242]
+ BL[243] BL[244] BL[245] BL[246] BL[247] BL[248] BL[249] BL[250] BL[251]
+ BL[252] BL[253] BL[254] BL[255] BLB[0] BLB[1] BLB[2] BLB[3] BLB[4] BLB[5]
+ BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15]
+ BLB[16] BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] BLB[24]
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] BLB[32] BLB[33]
+ BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] BLB[40] BLB[41] BLB[42]
+ BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] BLB[48] BLB[49] BLB[50] BLB[51]
+ BLB[52] BLB[53] BLB[54] BLB[55] BLB[56] BLB[57] BLB[58] BLB[59] BLB[60]
+ BLB[61] BLB[62] BLB[63] BLB[64] BLB[65] BLB[66] BLB[67] BLB[68] BLB[69]
+ BLB[70] BLB[71] BLB[72] BLB[73] BLB[74] BLB[75] BLB[76] BLB[77] BLB[78]
+ BLB[79] BLB[80] BLB[81] BLB[82] BLB[83] BLB[84] BLB[85] BLB[86] BLB[87]
+ BLB[88] BLB[89] BLB[90] BLB[91] BLB[92] BLB[93] BLB[94] BLB[95] BLB[96]
+ BLB[97] BLB[98] BLB[99] BLB[100] BLB[101] BLB[102] BLB[103] BLB[104] BLB[105]
+ BLB[106] BLB[107] BLB[108] BLB[109] BLB[110] BLB[111] BLB[112] BLB[113]
+ BLB[114] BLB[115] BLB[116] BLB[117] BLB[118] BLB[119] BLB[120] BLB[121]
+ BLB[122] BLB[123] BLB[124] BLB[125] BLB[126] BLB[127] BLB[128] BLB[129]
+ BLB[130] BLB[131] BLB[132] BLB[133] BLB[134] BLB[135] BLB[136] BLB[137]
+ BLB[138] BLB[139] BLB[140] BLB[141] BLB[142] BLB[143] BLB[144] BLB[145]
+ BLB[146] BLB[147] BLB[148] BLB[149] BLB[150] BLB[151] BLB[152] BLB[153]
+ BLB[154] BLB[155] BLB[156] BLB[157] BLB[158] BLB[159] BLB[160] BLB[161]
+ BLB[162] BLB[163] BLB[164] BLB[165] BLB[166] BLB[167] BLB[168] BLB[169]
+ BLB[170] BLB[171] BLB[172] BLB[173] BLB[174] BLB[175] BLB[176] BLB[177]
+ BLB[178] BLB[179] BLB[180] BLB[181] BLB[182] BLB[183] BLB[184] BLB[185]
+ BLB[186] BLB[187] BLB[188] BLB[189] BLB[190] BLB[191] BLB[192] BLB[193]
+ BLB[194] BLB[195] BLB[196] BLB[197] BLB[198] BLB[199] BLB[200] BLB[201]
+ BLB[202] BLB[203] BLB[204] BLB[205] BLB[206] BLB[207] BLB[208] BLB[209]
+ BLB[210] BLB[211] BLB[212] BLB[213] BLB[214] BLB[215] BLB[216] BLB[217]
+ BLB[218] BLB[219] BLB[220] BLB[221] BLB[222] BLB[223] BLB[224] BLB[225]
+ BLB[226] BLB[227] BLB[228] BLB[229] BLB[230] BLB[231] BLB[232] BLB[233]
+ BLB[234] BLB[235] BLB[236] BLB[237] BLB[238] BLB[239] BLB[240] BLB[241]
+ BLB[242] BLB[243] BLB[244] BLB[245] BLB[246] BLB[247] BLB[248] BLB[249]
+ BLB[250] BLB[251] BLB[252] BLB[253] BLB[254] BLB[255] WL[62] WL[63] VDDI VSSI
+ GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9] GBL[10]
+ GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18] GBL[19]
+ GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27] GBL[28]
+ GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36] GBL[37]
+ GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45] GBL[46]
+ GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54] GBL[55]
+ GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63] GBLB[0]
+ GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8] GBLB[9]
+ GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16] GBLB[17]
+ GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24] GBLB[25]
+ GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32] GBLB[33]
+ GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40] GBLB[41]
+ GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48] GBLB[49]
+ GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56] GBLB[57]
+ GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1] GW[2] GW[3]
+ GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15]
+ GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26]
+ GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37]
+ GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48]
+ GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59]
+ GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6]
+ GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16]
+ GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25]
+ GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34]
+ GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43]
+ GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52]
+ GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61]
+ GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_X
.ENDS

.SUBCKT S1AHSF400W40_LIO_MCB_F GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6]
+ GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16]
+ GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25]
+ GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34]
+ GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43]
+ GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52]
+ GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61]
+ GBL[62] GBL[63] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6]
+ GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15]
+ GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23]
+ GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31]
+ GBLB[32] GBLB[33] GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39]
+ GBLB[40] GBLB[41] GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47]
+ GBLB[48] GBLB[49] GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55]
+ GBLB[56] GBLB[57] GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] VDDHD
+ WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] WL[11]
+ WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] WL[22]
+ WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] WL[33]
+ WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] WL[44]
+ WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] WL[55]
+ WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] WL[64] WL[65] WL[66]
+ WL[67] WL[68] WL[69] WL[70] WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] WL[77]
+ WL[78] WL[79] WL[80] WL[81] WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] WL[88]
+ WL[89] WL[90] WL[91] WL[92] WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] WL[99]
+ WL[100] WL[101] WL[102] WL[103] WL[104] WL[105] WL[106] WL[107] WL[108]
+ WL[109] WL[110] WL[111] WL[112] WL[113] WL[114] WL[115] WL[116] WL[117]
+ WL[118] WL[119] WL[120] WL[121] WL[122] WL[123] WL[124] WL[125] WL[126]
+ WL[127] BLEQ_DN BLEQ_UP GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8]
+ GW[9] GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19]
+ GW[20] GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30]
+ GW[31] GW[32] GW[33] GW[34] GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41]
+ GW[42] GW[43] GW[44] GW[45] GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52]
+ GW[53] GW[54] GW[55] GW[56] GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63]
+ GWB[0] GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10]
+ GWB[11] GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19]
+ GWB[20] GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28]
+ GWB[29] GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37]
+ GWB[38] GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46]
+ GWB[47] GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55]
+ GWB[56] GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] RE SAEB WE
+ Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0]
+ Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] YL_LIO[0] YL_LIO[1]
+ VDDI VSSI
XCELL_ARR_DN_F BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] BL_DN[4] BL_DN[5] BL_DN[6]
+ BL_DN[7] BL_DN[8] BL_DN[9] BL_DN[10] BL_DN[11] BL_DN[12] BL_DN[13] BL_DN[14]
+ BL_DN[15] BL_DN[16] BL_DN[17] BL_DN[18] BL_DN[19] BL_DN[20] BL_DN[21]
+ BL_DN[22] BL_DN[23] BL_DN[24] BL_DN[25] BL_DN[26] BL_DN[27] BL_DN[28]
+ BL_DN[29] BL_DN[30] BL_DN[31] BL_DN[32] BL_DN[33] BL_DN[34] BL_DN[35]
+ BL_DN[36] BL_DN[37] BL_DN[38] BL_DN[39] BL_DN[40] BL_DN[41] BL_DN[42]
+ BL_DN[43] BL_DN[44] BL_DN[45] BL_DN[46] BL_DN[47] BL_DN[48] BL_DN[49]
+ BL_DN[50] BL_DN[51] BL_DN[52] BL_DN[53] BL_DN[54] BL_DN[55] BL_DN[56]
+ BL_DN[57] BL_DN[58] BL_DN[59] BL_DN[60] BL_DN[61] BL_DN[62] BL_DN[63]
+ BL_DN[64] BL_DN[65] BL_DN[66] BL_DN[67] BL_DN[68] BL_DN[69] BL_DN[70]
+ BL_DN[71] BL_DN[72] BL_DN[73] BL_DN[74] BL_DN[75] BL_DN[76] BL_DN[77]
+ BL_DN[78] BL_DN[79] BL_DN[80] BL_DN[81] BL_DN[82] BL_DN[83] BL_DN[84]
+ BL_DN[85] BL_DN[86] BL_DN[87] BL_DN[88] BL_DN[89] BL_DN[90] BL_DN[91]
+ BL_DN[92] BL_DN[93] BL_DN[94] BL_DN[95] BL_DN[96] BL_DN[97] BL_DN[98]
+ BL_DN[99] BL_DN[100] BL_DN[101] BL_DN[102] BL_DN[103] BL_DN[104] BL_DN[105]
+ BL_DN[106] BL_DN[107] BL_DN[108] BL_DN[109] BL_DN[110] BL_DN[111] BL_DN[112]
+ BL_DN[113] BL_DN[114] BL_DN[115] BL_DN[116] BL_DN[117] BL_DN[118] BL_DN[119]
+ BL_DN[120] BL_DN[121] BL_DN[122] BL_DN[123] BL_DN[124] BL_DN[125] BL_DN[126]
+ BL_DN[127] BL_DN[128] BL_DN[129] BL_DN[130] BL_DN[131] BL_DN[132] BL_DN[133]
+ BL_DN[134] BL_DN[135] BL_DN[136] BL_DN[137] BL_DN[138] BL_DN[139] BL_DN[140]
+ BL_DN[141] BL_DN[142] BL_DN[143] BL_DN[144] BL_DN[145] BL_DN[146] BL_DN[147]
+ BL_DN[148] BL_DN[149] BL_DN[150] BL_DN[151] BL_DN[152] BL_DN[153] BL_DN[154]
+ BL_DN[155] BL_DN[156] BL_DN[157] BL_DN[158] BL_DN[159] BL_DN[160] BL_DN[161]
+ BL_DN[162] BL_DN[163] BL_DN[164] BL_DN[165] BL_DN[166] BL_DN[167] BL_DN[168]
+ BL_DN[169] BL_DN[170] BL_DN[171] BL_DN[172] BL_DN[173] BL_DN[174] BL_DN[175]
+ BL_DN[176] BL_DN[177] BL_DN[178] BL_DN[179] BL_DN[180] BL_DN[181] BL_DN[182]
+ BL_DN[183] BL_DN[184] BL_DN[185] BL_DN[186] BL_DN[187] BL_DN[188] BL_DN[189]
+ BL_DN[190] BL_DN[191] BL_DN[192] BL_DN[193] BL_DN[194] BL_DN[195] BL_DN[196]
+ BL_DN[197] BL_DN[198] BL_DN[199] BL_DN[200] BL_DN[201] BL_DN[202] BL_DN[203]
+ BL_DN[204] BL_DN[205] BL_DN[206] BL_DN[207] BL_DN[208] BL_DN[209] BL_DN[210]
+ BL_DN[211] BL_DN[212] BL_DN[213] BL_DN[214] BL_DN[215] BL_DN[216] BL_DN[217]
+ BL_DN[218] BL_DN[219] BL_DN[220] BL_DN[221] BL_DN[222] BL_DN[223] BL_DN[224]
+ BL_DN[225] BL_DN[226] BL_DN[227] BL_DN[228] BL_DN[229] BL_DN[230] BL_DN[231]
+ BL_DN[232] BL_DN[233] BL_DN[234] BL_DN[235] BL_DN[236] BL_DN[237] BL_DN[238]
+ BL_DN[239] BL_DN[240] BL_DN[241] BL_DN[242] BL_DN[243] BL_DN[244] BL_DN[245]
+ BL_DN[246] BL_DN[247] BL_DN[248] BL_DN[249] BL_DN[250] BL_DN[251] BL_DN[252]
+ BL_DN[253] BL_DN[254] BL_DN[255] BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3]
+ BLB_DN[4] BLB_DN[5] BLB_DN[6] BLB_DN[7] BLB_DN[8] BLB_DN[9] BLB_DN[10]
+ BLB_DN[11] BLB_DN[12] BLB_DN[13] BLB_DN[14] BLB_DN[15] BLB_DN[16] BLB_DN[17]
+ BLB_DN[18] BLB_DN[19] BLB_DN[20] BLB_DN[21] BLB_DN[22] BLB_DN[23] BLB_DN[24]
+ BLB_DN[25] BLB_DN[26] BLB_DN[27] BLB_DN[28] BLB_DN[29] BLB_DN[30] BLB_DN[31]
+ BLB_DN[32] BLB_DN[33] BLB_DN[34] BLB_DN[35] BLB_DN[36] BLB_DN[37] BLB_DN[38]
+ BLB_DN[39] BLB_DN[40] BLB_DN[41] BLB_DN[42] BLB_DN[43] BLB_DN[44] BLB_DN[45]
+ BLB_DN[46] BLB_DN[47] BLB_DN[48] BLB_DN[49] BLB_DN[50] BLB_DN[51] BLB_DN[52]
+ BLB_DN[53] BLB_DN[54] BLB_DN[55] BLB_DN[56] BLB_DN[57] BLB_DN[58] BLB_DN[59]
+ BLB_DN[60] BLB_DN[61] BLB_DN[62] BLB_DN[63] BLB_DN[64] BLB_DN[65] BLB_DN[66]
+ BLB_DN[67] BLB_DN[68] BLB_DN[69] BLB_DN[70] BLB_DN[71] BLB_DN[72] BLB_DN[73]
+ BLB_DN[74] BLB_DN[75] BLB_DN[76] BLB_DN[77] BLB_DN[78] BLB_DN[79] BLB_DN[80]
+ BLB_DN[81] BLB_DN[82] BLB_DN[83] BLB_DN[84] BLB_DN[85] BLB_DN[86] BLB_DN[87]
+ BLB_DN[88] BLB_DN[89] BLB_DN[90] BLB_DN[91] BLB_DN[92] BLB_DN[93] BLB_DN[94]
+ BLB_DN[95] BLB_DN[96] BLB_DN[97] BLB_DN[98] BLB_DN[99] BLB_DN[100] BLB_DN[101]
+ BLB_DN[102] BLB_DN[103] BLB_DN[104] BLB_DN[105] BLB_DN[106] BLB_DN[107]
+ BLB_DN[108] BLB_DN[109] BLB_DN[110] BLB_DN[111] BLB_DN[112] BLB_DN[113]
+ BLB_DN[114] BLB_DN[115] BLB_DN[116] BLB_DN[117] BLB_DN[118] BLB_DN[119]
+ BLB_DN[120] BLB_DN[121] BLB_DN[122] BLB_DN[123] BLB_DN[124] BLB_DN[125]
+ BLB_DN[126] BLB_DN[127] BLB_DN[128] BLB_DN[129] BLB_DN[130] BLB_DN[131]
+ BLB_DN[132] BLB_DN[133] BLB_DN[134] BLB_DN[135] BLB_DN[136] BLB_DN[137]
+ BLB_DN[138] BLB_DN[139] BLB_DN[140] BLB_DN[141] BLB_DN[142] BLB_DN[143]
+ BLB_DN[144] BLB_DN[145] BLB_DN[146] BLB_DN[147] BLB_DN[148] BLB_DN[149]
+ BLB_DN[150] BLB_DN[151] BLB_DN[152] BLB_DN[153] BLB_DN[154] BLB_DN[155]
+ BLB_DN[156] BLB_DN[157] BLB_DN[158] BLB_DN[159] BLB_DN[160] BLB_DN[161]
+ BLB_DN[162] BLB_DN[163] BLB_DN[164] BLB_DN[165] BLB_DN[166] BLB_DN[167]
+ BLB_DN[168] BLB_DN[169] BLB_DN[170] BLB_DN[171] BLB_DN[172] BLB_DN[173]
+ BLB_DN[174] BLB_DN[175] BLB_DN[176] BLB_DN[177] BLB_DN[178] BLB_DN[179]
+ BLB_DN[180] BLB_DN[181] BLB_DN[182] BLB_DN[183] BLB_DN[184] BLB_DN[185]
+ BLB_DN[186] BLB_DN[187] BLB_DN[188] BLB_DN[189] BLB_DN[190] BLB_DN[191]
+ BLB_DN[192] BLB_DN[193] BLB_DN[194] BLB_DN[195] BLB_DN[196] BLB_DN[197]
+ BLB_DN[198] BLB_DN[199] BLB_DN[200] BLB_DN[201] BLB_DN[202] BLB_DN[203]
+ BLB_DN[204] BLB_DN[205] BLB_DN[206] BLB_DN[207] BLB_DN[208] BLB_DN[209]
+ BLB_DN[210] BLB_DN[211] BLB_DN[212] BLB_DN[213] BLB_DN[214] BLB_DN[215]
+ BLB_DN[216] BLB_DN[217] BLB_DN[218] BLB_DN[219] BLB_DN[220] BLB_DN[221]
+ BLB_DN[222] BLB_DN[223] BLB_DN[224] BLB_DN[225] BLB_DN[226] BLB_DN[227]
+ BLB_DN[228] BLB_DN[229] BLB_DN[230] BLB_DN[231] BLB_DN[232] BLB_DN[233]
+ BLB_DN[234] BLB_DN[235] BLB_DN[236] BLB_DN[237] BLB_DN[238] BLB_DN[239]
+ BLB_DN[240] BLB_DN[241] BLB_DN[242] BLB_DN[243] BLB_DN[244] BLB_DN[245]
+ BLB_DN[246] BLB_DN[247] BLB_DN[248] BLB_DN[249] BLB_DN[250] BLB_DN[251]
+ BLB_DN[252] BLB_DN[253] BLB_DN[254] BLB_DN[255] WL[0] WL[1] WL[2] WL[3] WL[4]
+ WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16]
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27]
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38]
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49]
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60]
+ WL[61] WL[62] WL[63] VDDI VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5]
+ GBL[6] GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15]
+ GBL[16] GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24]
+ GBL[25] GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33]
+ GBL[34] GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42]
+ GBL[43] GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51]
+ GBL[52] GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60]
+ GBL[61] GBL[62] GBL[63] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5]
+ GBLB[6] GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14]
+ GBLB[15] GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22]
+ GBLB[23] GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30]
+ GBLB[31] GBLB[32] GBLB[33] GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38]
+ GBLB[39] GBLB[40] GBLB[41] GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46]
+ GBLB[47] GBLB[48] GBLB[49] GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54]
+ GBLB[55] GBLB[56] GBLB[57] GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62]
+ GBLB[63] GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10]
+ GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21]
+ GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32]
+ GW[33] GW[34] GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43]
+ GW[44] GW[45] GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54]
+ GW[55] GW[56] GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1]
+ GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63]
+ S1AHSF400W40_CELL_ARR_XY_F
XCELL_ARR_UP_F BL_UP[0] BL_UP[1] BL_UP[2] BL_UP[3] BL_UP[4] BL_UP[5] BL_UP[6]
+ BL_UP[7] BL_UP[8] BL_UP[9] BL_UP[10] BL_UP[11] BL_UP[12] BL_UP[13] BL_UP[14]
+ BL_UP[15] BL_UP[16] BL_UP[17] BL_UP[18] BL_UP[19] BL_UP[20] BL_UP[21]
+ BL_UP[22] BL_UP[23] BL_UP[24] BL_UP[25] BL_UP[26] BL_UP[27] BL_UP[28]
+ BL_UP[29] BL_UP[30] BL_UP[31] BL_UP[32] BL_UP[33] BL_UP[34] BL_UP[35]
+ BL_UP[36] BL_UP[37] BL_UP[38] BL_UP[39] BL_UP[40] BL_UP[41] BL_UP[42]
+ BL_UP[43] BL_UP[44] BL_UP[45] BL_UP[46] BL_UP[47] BL_UP[48] BL_UP[49]
+ BL_UP[50] BL_UP[51] BL_UP[52] BL_UP[53] BL_UP[54] BL_UP[55] BL_UP[56]
+ BL_UP[57] BL_UP[58] BL_UP[59] BL_UP[60] BL_UP[61] BL_UP[62] BL_UP[63]
+ BL_UP[64] BL_UP[65] BL_UP[66] BL_UP[67] BL_UP[68] BL_UP[69] BL_UP[70]
+ BL_UP[71] BL_UP[72] BL_UP[73] BL_UP[74] BL_UP[75] BL_UP[76] BL_UP[77]
+ BL_UP[78] BL_UP[79] BL_UP[80] BL_UP[81] BL_UP[82] BL_UP[83] BL_UP[84]
+ BL_UP[85] BL_UP[86] BL_UP[87] BL_UP[88] BL_UP[89] BL_UP[90] BL_UP[91]
+ BL_UP[92] BL_UP[93] BL_UP[94] BL_UP[95] BL_UP[96] BL_UP[97] BL_UP[98]
+ BL_UP[99] BL_UP[100] BL_UP[101] BL_UP[102] BL_UP[103] BL_UP[104] BL_UP[105]
+ BL_UP[106] BL_UP[107] BL_UP[108] BL_UP[109] BL_UP[110] BL_UP[111] BL_UP[112]
+ BL_UP[113] BL_UP[114] BL_UP[115] BL_UP[116] BL_UP[117] BL_UP[118] BL_UP[119]
+ BL_UP[120] BL_UP[121] BL_UP[122] BL_UP[123] BL_UP[124] BL_UP[125] BL_UP[126]
+ BL_UP[127] BL_UP[128] BL_UP[129] BL_UP[130] BL_UP[131] BL_UP[132] BL_UP[133]
+ BL_UP[134] BL_UP[135] BL_UP[136] BL_UP[137] BL_UP[138] BL_UP[139] BL_UP[140]
+ BL_UP[141] BL_UP[142] BL_UP[143] BL_UP[144] BL_UP[145] BL_UP[146] BL_UP[147]
+ BL_UP[148] BL_UP[149] BL_UP[150] BL_UP[151] BL_UP[152] BL_UP[153] BL_UP[154]
+ BL_UP[155] BL_UP[156] BL_UP[157] BL_UP[158] BL_UP[159] BL_UP[160] BL_UP[161]
+ BL_UP[162] BL_UP[163] BL_UP[164] BL_UP[165] BL_UP[166] BL_UP[167] BL_UP[168]
+ BL_UP[169] BL_UP[170] BL_UP[171] BL_UP[172] BL_UP[173] BL_UP[174] BL_UP[175]
+ BL_UP[176] BL_UP[177] BL_UP[178] BL_UP[179] BL_UP[180] BL_UP[181] BL_UP[182]
+ BL_UP[183] BL_UP[184] BL_UP[185] BL_UP[186] BL_UP[187] BL_UP[188] BL_UP[189]
+ BL_UP[190] BL_UP[191] BL_UP[192] BL_UP[193] BL_UP[194] BL_UP[195] BL_UP[196]
+ BL_UP[197] BL_UP[198] BL_UP[199] BL_UP[200] BL_UP[201] BL_UP[202] BL_UP[203]
+ BL_UP[204] BL_UP[205] BL_UP[206] BL_UP[207] BL_UP[208] BL_UP[209] BL_UP[210]
+ BL_UP[211] BL_UP[212] BL_UP[213] BL_UP[214] BL_UP[215] BL_UP[216] BL_UP[217]
+ BL_UP[218] BL_UP[219] BL_UP[220] BL_UP[221] BL_UP[222] BL_UP[223] BL_UP[224]
+ BL_UP[225] BL_UP[226] BL_UP[227] BL_UP[228] BL_UP[229] BL_UP[230] BL_UP[231]
+ BL_UP[232] BL_UP[233] BL_UP[234] BL_UP[235] BL_UP[236] BL_UP[237] BL_UP[238]
+ BL_UP[239] BL_UP[240] BL_UP[241] BL_UP[242] BL_UP[243] BL_UP[244] BL_UP[245]
+ BL_UP[246] BL_UP[247] BL_UP[248] BL_UP[249] BL_UP[250] BL_UP[251] BL_UP[252]
+ BL_UP[253] BL_UP[254] BL_UP[255] BLB_UP[0] BLB_UP[1] BLB_UP[2] BLB_UP[3]
+ BLB_UP[4] BLB_UP[5] BLB_UP[6] BLB_UP[7] BLB_UP[8] BLB_UP[9] BLB_UP[10]
+ BLB_UP[11] BLB_UP[12] BLB_UP[13] BLB_UP[14] BLB_UP[15] BLB_UP[16] BLB_UP[17]
+ BLB_UP[18] BLB_UP[19] BLB_UP[20] BLB_UP[21] BLB_UP[22] BLB_UP[23] BLB_UP[24]
+ BLB_UP[25] BLB_UP[26] BLB_UP[27] BLB_UP[28] BLB_UP[29] BLB_UP[30] BLB_UP[31]
+ BLB_UP[32] BLB_UP[33] BLB_UP[34] BLB_UP[35] BLB_UP[36] BLB_UP[37] BLB_UP[38]
+ BLB_UP[39] BLB_UP[40] BLB_UP[41] BLB_UP[42] BLB_UP[43] BLB_UP[44] BLB_UP[45]
+ BLB_UP[46] BLB_UP[47] BLB_UP[48] BLB_UP[49] BLB_UP[50] BLB_UP[51] BLB_UP[52]
+ BLB_UP[53] BLB_UP[54] BLB_UP[55] BLB_UP[56] BLB_UP[57] BLB_UP[58] BLB_UP[59]
+ BLB_UP[60] BLB_UP[61] BLB_UP[62] BLB_UP[63] BLB_UP[64] BLB_UP[65] BLB_UP[66]
+ BLB_UP[67] BLB_UP[68] BLB_UP[69] BLB_UP[70] BLB_UP[71] BLB_UP[72] BLB_UP[73]
+ BLB_UP[74] BLB_UP[75] BLB_UP[76] BLB_UP[77] BLB_UP[78] BLB_UP[79] BLB_UP[80]
+ BLB_UP[81] BLB_UP[82] BLB_UP[83] BLB_UP[84] BLB_UP[85] BLB_UP[86] BLB_UP[87]
+ BLB_UP[88] BLB_UP[89] BLB_UP[90] BLB_UP[91] BLB_UP[92] BLB_UP[93] BLB_UP[94]
+ BLB_UP[95] BLB_UP[96] BLB_UP[97] BLB_UP[98] BLB_UP[99] BLB_UP[100] BLB_UP[101]
+ BLB_UP[102] BLB_UP[103] BLB_UP[104] BLB_UP[105] BLB_UP[106] BLB_UP[107]
+ BLB_UP[108] BLB_UP[109] BLB_UP[110] BLB_UP[111] BLB_UP[112] BLB_UP[113]
+ BLB_UP[114] BLB_UP[115] BLB_UP[116] BLB_UP[117] BLB_UP[118] BLB_UP[119]
+ BLB_UP[120] BLB_UP[121] BLB_UP[122] BLB_UP[123] BLB_UP[124] BLB_UP[125]
+ BLB_UP[126] BLB_UP[127] BLB_UP[128] BLB_UP[129] BLB_UP[130] BLB_UP[131]
+ BLB_UP[132] BLB_UP[133] BLB_UP[134] BLB_UP[135] BLB_UP[136] BLB_UP[137]
+ BLB_UP[138] BLB_UP[139] BLB_UP[140] BLB_UP[141] BLB_UP[142] BLB_UP[143]
+ BLB_UP[144] BLB_UP[145] BLB_UP[146] BLB_UP[147] BLB_UP[148] BLB_UP[149]
+ BLB_UP[150] BLB_UP[151] BLB_UP[152] BLB_UP[153] BLB_UP[154] BLB_UP[155]
+ BLB_UP[156] BLB_UP[157] BLB_UP[158] BLB_UP[159] BLB_UP[160] BLB_UP[161]
+ BLB_UP[162] BLB_UP[163] BLB_UP[164] BLB_UP[165] BLB_UP[166] BLB_UP[167]
+ BLB_UP[168] BLB_UP[169] BLB_UP[170] BLB_UP[171] BLB_UP[172] BLB_UP[173]
+ BLB_UP[174] BLB_UP[175] BLB_UP[176] BLB_UP[177] BLB_UP[178] BLB_UP[179]
+ BLB_UP[180] BLB_UP[181] BLB_UP[182] BLB_UP[183] BLB_UP[184] BLB_UP[185]
+ BLB_UP[186] BLB_UP[187] BLB_UP[188] BLB_UP[189] BLB_UP[190] BLB_UP[191]
+ BLB_UP[192] BLB_UP[193] BLB_UP[194] BLB_UP[195] BLB_UP[196] BLB_UP[197]
+ BLB_UP[198] BLB_UP[199] BLB_UP[200] BLB_UP[201] BLB_UP[202] BLB_UP[203]
+ BLB_UP[204] BLB_UP[205] BLB_UP[206] BLB_UP[207] BLB_UP[208] BLB_UP[209]
+ BLB_UP[210] BLB_UP[211] BLB_UP[212] BLB_UP[213] BLB_UP[214] BLB_UP[215]
+ BLB_UP[216] BLB_UP[217] BLB_UP[218] BLB_UP[219] BLB_UP[220] BLB_UP[221]
+ BLB_UP[222] BLB_UP[223] BLB_UP[224] BLB_UP[225] BLB_UP[226] BLB_UP[227]
+ BLB_UP[228] BLB_UP[229] BLB_UP[230] BLB_UP[231] BLB_UP[232] BLB_UP[233]
+ BLB_UP[234] BLB_UP[235] BLB_UP[236] BLB_UP[237] BLB_UP[238] BLB_UP[239]
+ BLB_UP[240] BLB_UP[241] BLB_UP[242] BLB_UP[243] BLB_UP[244] BLB_UP[245]
+ BLB_UP[246] BLB_UP[247] BLB_UP[248] BLB_UP[249] BLB_UP[250] BLB_UP[251]
+ BLB_UP[252] BLB_UP[253] BLB_UP[254] BLB_UP[255] WL[64] WL[65] WL[66] WL[67]
+ WL[68] WL[69] WL[70] WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78]
+ WL[79] WL[80] WL[81] WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89]
+ WL[90] WL[91] WL[92] WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100]
+ WL[101] WL[102] WL[103] WL[104] WL[105] WL[106] WL[107] WL[108] WL[109]
+ WL[110] WL[111] WL[112] WL[113] WL[114] WL[115] WL[116] WL[117] WL[118]
+ WL[119] WL[120] WL[121] WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] VDDI
+ VSSI GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9]
+ GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18]
+ GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27]
+ GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36]
+ GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45]
+ GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54]
+ GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63]
+ GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8]
+ GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16]
+ GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24]
+ GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32]
+ GBLB[33] GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40]
+ GBLB[41] GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48]
+ GBLB[49] GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56]
+ GBLB[57] GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1]
+ GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13]
+ GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24]
+ GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35]
+ GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46]
+ GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57]
+ GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4]
+ GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14]
+ GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23]
+ GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32]
+ GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41]
+ GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50]
+ GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59]
+ GWB[60] GWB[61] GWB[62] GWB[63] S1AHSF400W40_CELL_ARR_XY_F
XLIO_M4_0 BLB_DN[0] BLB_DN[1] BLB_DN[2] BLB_DN[3] BLB_UP[0] BLB_UP[1] BLB_UP[2]
+ BLB_UP[3] BLEQ_DN BLEQ_UP BL_DN[0] BL_DN[1] BL_DN[2] BL_DN[3] BL_UP[0]
+ BL_UP[1] BL_UP[2] BL_UP[3] GBL[0] GBLB[0] GW[0] GWB[0] RE SAEB VDDHD VDDI VSSI
+ WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6]
+ Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ S1AHSF400W40_LIO_M4
XLIO_M4_1 BLB_DN[4] BLB_DN[5] BLB_DN[6] BLB_DN[7] BLB_UP[4] BLB_UP[5] BLB_UP[6]
+ BLB_UP[7] BLEQ_DN BLEQ_UP BL_DN[4] BL_DN[5] BL_DN[6] BL_DN[7] BL_UP[4]
+ BL_UP[5] BL_UP[6] BL_UP[7] GBL[1] GBLB[1] GW[1] GWB[1] RE SAEB VDDHD VDDI VSSI
+ WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6]
+ Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7]
+ S1AHSF400W40_LIO_M4
XLIO_M4_2 BLB_DN[8] BLB_DN[9] BLB_DN[10] BLB_DN[11] BLB_UP[8] BLB_UP[9]
+ BLB_UP[10] BLB_UP[11] BLEQ_DN BLEQ_UP BL_DN[8] BL_DN[9] BL_DN[10] BL_DN[11]
+ BL_UP[8] BL_UP[9] BL_UP[10] BL_UP[11] GBL[2] GBLB[2] GW[2] GWB[2] RE SAEB
+ VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4]
+ Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5]
+ Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_3 BLB_DN[12] BLB_DN[13] BLB_DN[14] BLB_DN[15] BLB_UP[12] BLB_UP[13]
+ BLB_UP[14] BLB_UP[15] BLEQ_DN BLEQ_UP BL_DN[12] BL_DN[13] BL_DN[14] BL_DN[15]
+ BL_UP[12] BL_UP[13] BL_UP[14] BL_UP[15] GBL[3] GBLB[3] GW[3] GWB[3] RE SAEB
+ VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4]
+ Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5]
+ Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_4 BLB_DN[16] BLB_DN[17] BLB_DN[18] BLB_DN[19] BLB_UP[16] BLB_UP[17]
+ BLB_UP[18] BLB_UP[19] BLEQ_DN BLEQ_UP BL_DN[16] BL_DN[17] BL_DN[18] BL_DN[19]
+ BL_UP[16] BL_UP[17] BL_UP[18] BL_UP[19] GBL[4] GBLB[4] GW[4] GWB[4] RE SAEB
+ VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4]
+ Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5]
+ Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_5 BLB_DN[20] BLB_DN[21] BLB_DN[22] BLB_DN[23] BLB_UP[20] BLB_UP[21]
+ BLB_UP[22] BLB_UP[23] BLEQ_DN BLEQ_UP BL_DN[20] BL_DN[21] BL_DN[22] BL_DN[23]
+ BL_UP[20] BL_UP[21] BL_UP[22] BL_UP[23] GBL[5] GBLB[5] GW[5] GWB[5] RE SAEB
+ VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4]
+ Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5]
+ Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_6 BLB_DN[24] BLB_DN[25] BLB_DN[26] BLB_DN[27] BLB_UP[24] BLB_UP[25]
+ BLB_UP[26] BLB_UP[27] BLEQ_DN BLEQ_UP BL_DN[24] BL_DN[25] BL_DN[26] BL_DN[27]
+ BL_UP[24] BL_UP[25] BL_UP[26] BL_UP[27] GBL[6] GBLB[6] GW[6] GWB[6] RE SAEB
+ VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4]
+ Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5]
+ Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_7 BLB_DN[28] BLB_DN[29] BLB_DN[30] BLB_DN[31] BLB_UP[28] BLB_UP[29]
+ BLB_UP[30] BLB_UP[31] BLEQ_DN BLEQ_UP BL_DN[28] BL_DN[29] BL_DN[30] BL_DN[31]
+ BL_UP[28] BL_UP[29] BL_UP[30] BL_UP[31] GBL[7] GBLB[7] GW[7] GWB[7] RE SAEB
+ VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4]
+ Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5]
+ Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_8 BLB_DN[32] BLB_DN[33] BLB_DN[34] BLB_DN[35] BLB_UP[32] BLB_UP[33]
+ BLB_UP[34] BLB_UP[35] BLEQ_DN BLEQ_UP BL_DN[32] BL_DN[33] BL_DN[34] BL_DN[35]
+ BL_UP[32] BL_UP[33] BL_UP[34] BL_UP[35] GBL[8] GBLB[8] GW[8] GWB[8] RE SAEB
+ VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4]
+ Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5]
+ Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_9 BLB_DN[36] BLB_DN[37] BLB_DN[38] BLB_DN[39] BLB_UP[36] BLB_UP[37]
+ BLB_UP[38] BLB_UP[39] BLEQ_DN BLEQ_UP BL_DN[36] BL_DN[37] BL_DN[38] BL_DN[39]
+ BL_UP[36] BL_UP[37] BL_UP[38] BL_UP[39] GBL[9] GBLB[9] GW[9] GWB[9] RE SAEB
+ VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4]
+ Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5]
+ Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_10 BLB_DN[40] BLB_DN[41] BLB_DN[42] BLB_DN[43] BLB_UP[40] BLB_UP[41]
+ BLB_UP[42] BLB_UP[43] BLEQ_DN BLEQ_UP BL_DN[40] BL_DN[41] BL_DN[42] BL_DN[43]
+ BL_UP[40] BL_UP[41] BL_UP[42] BL_UP[43] GBL[10] GBLB[10] GW[10] GWB[10] RE
+ SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_11 BLB_DN[44] BLB_DN[45] BLB_DN[46] BLB_DN[47] BLB_UP[44] BLB_UP[45]
+ BLB_UP[46] BLB_UP[47] BLEQ_DN BLEQ_UP BL_DN[44] BL_DN[45] BL_DN[46] BL_DN[47]
+ BL_UP[44] BL_UP[45] BL_UP[46] BL_UP[47] GBL[11] GBLB[11] GW[11] GWB[11] RE
+ SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_12 BLB_DN[48] BLB_DN[49] BLB_DN[50] BLB_DN[51] BLB_UP[48] BLB_UP[49]
+ BLB_UP[50] BLB_UP[51] BLEQ_DN BLEQ_UP BL_DN[48] BL_DN[49] BL_DN[50] BL_DN[51]
+ BL_UP[48] BL_UP[49] BL_UP[50] BL_UP[51] GBL[12] GBLB[12] GW[12] GWB[12] RE
+ SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_13 BLB_DN[52] BLB_DN[53] BLB_DN[54] BLB_DN[55] BLB_UP[52] BLB_UP[53]
+ BLB_UP[54] BLB_UP[55] BLEQ_DN BLEQ_UP BL_DN[52] BL_DN[53] BL_DN[54] BL_DN[55]
+ BL_UP[52] BL_UP[53] BL_UP[54] BL_UP[55] GBL[13] GBLB[13] GW[13] GWB[13] RE
+ SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_14 BLB_DN[56] BLB_DN[57] BLB_DN[58] BLB_DN[59] BLB_UP[56] BLB_UP[57]
+ BLB_UP[58] BLB_UP[59] BLEQ_DN BLEQ_UP BL_DN[56] BL_DN[57] BL_DN[58] BL_DN[59]
+ BL_UP[56] BL_UP[57] BL_UP[58] BL_UP[59] GBL[14] GBLB[14] GW[14] GWB[14] RE
+ SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_15 BLB_DN[60] BLB_DN[61] BLB_DN[62] BLB_DN[63] BLB_UP[60] BLB_UP[61]
+ BLB_UP[62] BLB_UP[63] BLEQ_DN BLEQ_UP BL_DN[60] BL_DN[61] BL_DN[62] BL_DN[63]
+ BL_UP[60] BL_UP[61] BL_UP[62] BL_UP[63] GBL[15] GBLB[15] GW[15] GWB[15] RE
+ SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_16 BLB_DN[64] BLB_DN[65] BLB_DN[66] BLB_DN[67] BLB_UP[64] BLB_UP[65]
+ BLB_UP[66] BLB_UP[67] BLEQ_DN BLEQ_UP BL_DN[64] BL_DN[65] BL_DN[66] BL_DN[67]
+ BL_UP[64] BL_UP[65] BL_UP[66] BL_UP[67] GBL[16] GBLB[16] GW[16] GWB[16] RE
+ SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_17 BLB_DN[68] BLB_DN[69] BLB_DN[70] BLB_DN[71] BLB_UP[68] BLB_UP[69]
+ BLB_UP[70] BLB_UP[71] BLEQ_DN BLEQ_UP BL_DN[68] BL_DN[69] BL_DN[70] BL_DN[71]
+ BL_UP[68] BL_UP[69] BL_UP[70] BL_UP[71] GBL[17] GBLB[17] GW[17] GWB[17] RE
+ SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_18 BLB_DN[72] BLB_DN[73] BLB_DN[74] BLB_DN[75] BLB_UP[72] BLB_UP[73]
+ BLB_UP[74] BLB_UP[75] BLEQ_DN BLEQ_UP BL_DN[72] BL_DN[73] BL_DN[74] BL_DN[75]
+ BL_UP[72] BL_UP[73] BL_UP[74] BL_UP[75] GBL[18] GBLB[18] GW[18] GWB[18] RE
+ SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_19 BLB_DN[76] BLB_DN[77] BLB_DN[78] BLB_DN[79] BLB_UP[76] BLB_UP[77]
+ BLB_UP[78] BLB_UP[79] BLEQ_DN BLEQ_UP BL_DN[76] BL_DN[77] BL_DN[78] BL_DN[79]
+ BL_UP[76] BL_UP[77] BL_UP[78] BL_UP[79] GBL[19] GBLB[19] GW[19] GWB[19] RE
+ SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_20 BLB_DN[80] BLB_DN[81] BLB_DN[82] BLB_DN[83] BLB_UP[80] BLB_UP[81]
+ BLB_UP[82] BLB_UP[83] BLEQ_DN BLEQ_UP BL_DN[80] BL_DN[81] BL_DN[82] BL_DN[83]
+ BL_UP[80] BL_UP[81] BL_UP[82] BL_UP[83] GBL[20] GBLB[20] GW[20] GWB[20] RE
+ SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_21 BLB_DN[84] BLB_DN[85] BLB_DN[86] BLB_DN[87] BLB_UP[84] BLB_UP[85]
+ BLB_UP[86] BLB_UP[87] BLEQ_DN BLEQ_UP BL_DN[84] BL_DN[85] BL_DN[86] BL_DN[87]
+ BL_UP[84] BL_UP[85] BL_UP[86] BL_UP[87] GBL[21] GBLB[21] GW[21] GWB[21] RE
+ SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_22 BLB_DN[88] BLB_DN[89] BLB_DN[90] BLB_DN[91] BLB_UP[88] BLB_UP[89]
+ BLB_UP[90] BLB_UP[91] BLEQ_DN BLEQ_UP BL_DN[88] BL_DN[89] BL_DN[90] BL_DN[91]
+ BL_UP[88] BL_UP[89] BL_UP[90] BL_UP[91] GBL[22] GBLB[22] GW[22] GWB[22] RE
+ SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_23 BLB_DN[92] BLB_DN[93] BLB_DN[94] BLB_DN[95] BLB_UP[92] BLB_UP[93]
+ BLB_UP[94] BLB_UP[95] BLEQ_DN BLEQ_UP BL_DN[92] BL_DN[93] BL_DN[94] BL_DN[95]
+ BL_UP[92] BL_UP[93] BL_UP[94] BL_UP[95] GBL[23] GBLB[23] GW[23] GWB[23] RE
+ SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_24 BLB_DN[96] BLB_DN[97] BLB_DN[98] BLB_DN[99] BLB_UP[96] BLB_UP[97]
+ BLB_UP[98] BLB_UP[99] BLEQ_DN BLEQ_UP BL_DN[96] BL_DN[97] BL_DN[98] BL_DN[99]
+ BL_UP[96] BL_UP[97] BL_UP[98] BL_UP[99] GBL[24] GBLB[24] GW[24] GWB[24] RE
+ SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0] Y_DN[1] Y_DN[2] Y_DN[3]
+ Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1] Y_UP[2] Y_UP[3] Y_UP[4]
+ Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_25 BLB_DN[100] BLB_DN[101] BLB_DN[102] BLB_DN[103] BLB_UP[100]
+ BLB_UP[101] BLB_UP[102] BLB_UP[103] BLEQ_DN BLEQ_UP BL_DN[100] BL_DN[101]
+ BL_DN[102] BL_DN[103] BL_UP[100] BL_UP[101] BL_UP[102] BL_UP[103] GBL[25]
+ GBLB[25] GW[25] GWB[25] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_26 BLB_DN[104] BLB_DN[105] BLB_DN[106] BLB_DN[107] BLB_UP[104]
+ BLB_UP[105] BLB_UP[106] BLB_UP[107] BLEQ_DN BLEQ_UP BL_DN[104] BL_DN[105]
+ BL_DN[106] BL_DN[107] BL_UP[104] BL_UP[105] BL_UP[106] BL_UP[107] GBL[26]
+ GBLB[26] GW[26] GWB[26] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_27 BLB_DN[108] BLB_DN[109] BLB_DN[110] BLB_DN[111] BLB_UP[108]
+ BLB_UP[109] BLB_UP[110] BLB_UP[111] BLEQ_DN BLEQ_UP BL_DN[108] BL_DN[109]
+ BL_DN[110] BL_DN[111] BL_UP[108] BL_UP[109] BL_UP[110] BL_UP[111] GBL[27]
+ GBLB[27] GW[27] GWB[27] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_28 BLB_DN[112] BLB_DN[113] BLB_DN[114] BLB_DN[115] BLB_UP[112]
+ BLB_UP[113] BLB_UP[114] BLB_UP[115] BLEQ_DN BLEQ_UP BL_DN[112] BL_DN[113]
+ BL_DN[114] BL_DN[115] BL_UP[112] BL_UP[113] BL_UP[114] BL_UP[115] GBL[28]
+ GBLB[28] GW[28] GWB[28] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_29 BLB_DN[116] BLB_DN[117] BLB_DN[118] BLB_DN[119] BLB_UP[116]
+ BLB_UP[117] BLB_UP[118] BLB_UP[119] BLEQ_DN BLEQ_UP BL_DN[116] BL_DN[117]
+ BL_DN[118] BL_DN[119] BL_UP[116] BL_UP[117] BL_UP[118] BL_UP[119] GBL[29]
+ GBLB[29] GW[29] GWB[29] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_30 BLB_DN[120] BLB_DN[121] BLB_DN[122] BLB_DN[123] BLB_UP[120]
+ BLB_UP[121] BLB_UP[122] BLB_UP[123] BLEQ_DN BLEQ_UP BL_DN[120] BL_DN[121]
+ BL_DN[122] BL_DN[123] BL_UP[120] BL_UP[121] BL_UP[122] BL_UP[123] GBL[30]
+ GBLB[30] GW[30] GWB[30] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_31 BLB_DN[124] BLB_DN[125] BLB_DN[126] BLB_DN[127] BLB_UP[124]
+ BLB_UP[125] BLB_UP[126] BLB_UP[127] BLEQ_DN BLEQ_UP BL_DN[124] BL_DN[125]
+ BL_DN[126] BL_DN[127] BL_UP[124] BL_UP[125] BL_UP[126] BL_UP[127] GBL[31]
+ GBLB[31] GW[31] GWB[31] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_32 BLB_DN[128] BLB_DN[129] BLB_DN[130] BLB_DN[131] BLB_UP[128]
+ BLB_UP[129] BLB_UP[130] BLB_UP[131] BLEQ_DN BLEQ_UP BL_DN[128] BL_DN[129]
+ BL_DN[130] BL_DN[131] BL_UP[128] BL_UP[129] BL_UP[130] BL_UP[131] GBL[32]
+ GBLB[32] GW[32] GWB[32] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_33 BLB_DN[132] BLB_DN[133] BLB_DN[134] BLB_DN[135] BLB_UP[132]
+ BLB_UP[133] BLB_UP[134] BLB_UP[135] BLEQ_DN BLEQ_UP BL_DN[132] BL_DN[133]
+ BL_DN[134] BL_DN[135] BL_UP[132] BL_UP[133] BL_UP[134] BL_UP[135] GBL[33]
+ GBLB[33] GW[33] GWB[33] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_34 BLB_DN[136] BLB_DN[137] BLB_DN[138] BLB_DN[139] BLB_UP[136]
+ BLB_UP[137] BLB_UP[138] BLB_UP[139] BLEQ_DN BLEQ_UP BL_DN[136] BL_DN[137]
+ BL_DN[138] BL_DN[139] BL_UP[136] BL_UP[137] BL_UP[138] BL_UP[139] GBL[34]
+ GBLB[34] GW[34] GWB[34] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_35 BLB_DN[140] BLB_DN[141] BLB_DN[142] BLB_DN[143] BLB_UP[140]
+ BLB_UP[141] BLB_UP[142] BLB_UP[143] BLEQ_DN BLEQ_UP BL_DN[140] BL_DN[141]
+ BL_DN[142] BL_DN[143] BL_UP[140] BL_UP[141] BL_UP[142] BL_UP[143] GBL[35]
+ GBLB[35] GW[35] GWB[35] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_36 BLB_DN[144] BLB_DN[145] BLB_DN[146] BLB_DN[147] BLB_UP[144]
+ BLB_UP[145] BLB_UP[146] BLB_UP[147] BLEQ_DN BLEQ_UP BL_DN[144] BL_DN[145]
+ BL_DN[146] BL_DN[147] BL_UP[144] BL_UP[145] BL_UP[146] BL_UP[147] GBL[36]
+ GBLB[36] GW[36] GWB[36] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_37 BLB_DN[148] BLB_DN[149] BLB_DN[150] BLB_DN[151] BLB_UP[148]
+ BLB_UP[149] BLB_UP[150] BLB_UP[151] BLEQ_DN BLEQ_UP BL_DN[148] BL_DN[149]
+ BL_DN[150] BL_DN[151] BL_UP[148] BL_UP[149] BL_UP[150] BL_UP[151] GBL[37]
+ GBLB[37] GW[37] GWB[37] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_38 BLB_DN[152] BLB_DN[153] BLB_DN[154] BLB_DN[155] BLB_UP[152]
+ BLB_UP[153] BLB_UP[154] BLB_UP[155] BLEQ_DN BLEQ_UP BL_DN[152] BL_DN[153]
+ BL_DN[154] BL_DN[155] BL_UP[152] BL_UP[153] BL_UP[154] BL_UP[155] GBL[38]
+ GBLB[38] GW[38] GWB[38] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_39 BLB_DN[156] BLB_DN[157] BLB_DN[158] BLB_DN[159] BLB_UP[156]
+ BLB_UP[157] BLB_UP[158] BLB_UP[159] BLEQ_DN BLEQ_UP BL_DN[156] BL_DN[157]
+ BL_DN[158] BL_DN[159] BL_UP[156] BL_UP[157] BL_UP[158] BL_UP[159] GBL[39]
+ GBLB[39] GW[39] GWB[39] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_40 BLB_DN[160] BLB_DN[161] BLB_DN[162] BLB_DN[163] BLB_UP[160]
+ BLB_UP[161] BLB_UP[162] BLB_UP[163] BLEQ_DN BLEQ_UP BL_DN[160] BL_DN[161]
+ BL_DN[162] BL_DN[163] BL_UP[160] BL_UP[161] BL_UP[162] BL_UP[163] GBL[40]
+ GBLB[40] GW[40] GWB[40] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_41 BLB_DN[164] BLB_DN[165] BLB_DN[166] BLB_DN[167] BLB_UP[164]
+ BLB_UP[165] BLB_UP[166] BLB_UP[167] BLEQ_DN BLEQ_UP BL_DN[164] BL_DN[165]
+ BL_DN[166] BL_DN[167] BL_UP[164] BL_UP[165] BL_UP[166] BL_UP[167] GBL[41]
+ GBLB[41] GW[41] GWB[41] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_42 BLB_DN[168] BLB_DN[169] BLB_DN[170] BLB_DN[171] BLB_UP[168]
+ BLB_UP[169] BLB_UP[170] BLB_UP[171] BLEQ_DN BLEQ_UP BL_DN[168] BL_DN[169]
+ BL_DN[170] BL_DN[171] BL_UP[168] BL_UP[169] BL_UP[170] BL_UP[171] GBL[42]
+ GBLB[42] GW[42] GWB[42] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_43 BLB_DN[172] BLB_DN[173] BLB_DN[174] BLB_DN[175] BLB_UP[172]
+ BLB_UP[173] BLB_UP[174] BLB_UP[175] BLEQ_DN BLEQ_UP BL_DN[172] BL_DN[173]
+ BL_DN[174] BL_DN[175] BL_UP[172] BL_UP[173] BL_UP[174] BL_UP[175] GBL[43]
+ GBLB[43] GW[43] GWB[43] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_44 BLB_DN[176] BLB_DN[177] BLB_DN[178] BLB_DN[179] BLB_UP[176]
+ BLB_UP[177] BLB_UP[178] BLB_UP[179] BLEQ_DN BLEQ_UP BL_DN[176] BL_DN[177]
+ BL_DN[178] BL_DN[179] BL_UP[176] BL_UP[177] BL_UP[178] BL_UP[179] GBL[44]
+ GBLB[44] GW[44] GWB[44] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_45 BLB_DN[180] BLB_DN[181] BLB_DN[182] BLB_DN[183] BLB_UP[180]
+ BLB_UP[181] BLB_UP[182] BLB_UP[183] BLEQ_DN BLEQ_UP BL_DN[180] BL_DN[181]
+ BL_DN[182] BL_DN[183] BL_UP[180] BL_UP[181] BL_UP[182] BL_UP[183] GBL[45]
+ GBLB[45] GW[45] GWB[45] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_46 BLB_DN[184] BLB_DN[185] BLB_DN[186] BLB_DN[187] BLB_UP[184]
+ BLB_UP[185] BLB_UP[186] BLB_UP[187] BLEQ_DN BLEQ_UP BL_DN[184] BL_DN[185]
+ BL_DN[186] BL_DN[187] BL_UP[184] BL_UP[185] BL_UP[186] BL_UP[187] GBL[46]
+ GBLB[46] GW[46] GWB[46] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_47 BLB_DN[188] BLB_DN[189] BLB_DN[190] BLB_DN[191] BLB_UP[188]
+ BLB_UP[189] BLB_UP[190] BLB_UP[191] BLEQ_DN BLEQ_UP BL_DN[188] BL_DN[189]
+ BL_DN[190] BL_DN[191] BL_UP[188] BL_UP[189] BL_UP[190] BL_UP[191] GBL[47]
+ GBLB[47] GW[47] GWB[47] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_48 BLB_DN[192] BLB_DN[193] BLB_DN[194] BLB_DN[195] BLB_UP[192]
+ BLB_UP[193] BLB_UP[194] BLB_UP[195] BLEQ_DN BLEQ_UP BL_DN[192] BL_DN[193]
+ BL_DN[194] BL_DN[195] BL_UP[192] BL_UP[193] BL_UP[194] BL_UP[195] GBL[48]
+ GBLB[48] GW[48] GWB[48] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_49 BLB_DN[196] BLB_DN[197] BLB_DN[198] BLB_DN[199] BLB_UP[196]
+ BLB_UP[197] BLB_UP[198] BLB_UP[199] BLEQ_DN BLEQ_UP BL_DN[196] BL_DN[197]
+ BL_DN[198] BL_DN[199] BL_UP[196] BL_UP[197] BL_UP[198] BL_UP[199] GBL[49]
+ GBLB[49] GW[49] GWB[49] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_50 BLB_DN[200] BLB_DN[201] BLB_DN[202] BLB_DN[203] BLB_UP[200]
+ BLB_UP[201] BLB_UP[202] BLB_UP[203] BLEQ_DN BLEQ_UP BL_DN[200] BL_DN[201]
+ BL_DN[202] BL_DN[203] BL_UP[200] BL_UP[201] BL_UP[202] BL_UP[203] GBL[50]
+ GBLB[50] GW[50] GWB[50] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_51 BLB_DN[204] BLB_DN[205] BLB_DN[206] BLB_DN[207] BLB_UP[204]
+ BLB_UP[205] BLB_UP[206] BLB_UP[207] BLEQ_DN BLEQ_UP BL_DN[204] BL_DN[205]
+ BL_DN[206] BL_DN[207] BL_UP[204] BL_UP[205] BL_UP[206] BL_UP[207] GBL[51]
+ GBLB[51] GW[51] GWB[51] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_52 BLB_DN[208] BLB_DN[209] BLB_DN[210] BLB_DN[211] BLB_UP[208]
+ BLB_UP[209] BLB_UP[210] BLB_UP[211] BLEQ_DN BLEQ_UP BL_DN[208] BL_DN[209]
+ BL_DN[210] BL_DN[211] BL_UP[208] BL_UP[209] BL_UP[210] BL_UP[211] GBL[52]
+ GBLB[52] GW[52] GWB[52] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_53 BLB_DN[212] BLB_DN[213] BLB_DN[214] BLB_DN[215] BLB_UP[212]
+ BLB_UP[213] BLB_UP[214] BLB_UP[215] BLEQ_DN BLEQ_UP BL_DN[212] BL_DN[213]
+ BL_DN[214] BL_DN[215] BL_UP[212] BL_UP[213] BL_UP[214] BL_UP[215] GBL[53]
+ GBLB[53] GW[53] GWB[53] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_54 BLB_DN[216] BLB_DN[217] BLB_DN[218] BLB_DN[219] BLB_UP[216]
+ BLB_UP[217] BLB_UP[218] BLB_UP[219] BLEQ_DN BLEQ_UP BL_DN[216] BL_DN[217]
+ BL_DN[218] BL_DN[219] BL_UP[216] BL_UP[217] BL_UP[218] BL_UP[219] GBL[54]
+ GBLB[54] GW[54] GWB[54] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_55 BLB_DN[220] BLB_DN[221] BLB_DN[222] BLB_DN[223] BLB_UP[220]
+ BLB_UP[221] BLB_UP[222] BLB_UP[223] BLEQ_DN BLEQ_UP BL_DN[220] BL_DN[221]
+ BL_DN[222] BL_DN[223] BL_UP[220] BL_UP[221] BL_UP[222] BL_UP[223] GBL[55]
+ GBLB[55] GW[55] GWB[55] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_56 BLB_DN[224] BLB_DN[225] BLB_DN[226] BLB_DN[227] BLB_UP[224]
+ BLB_UP[225] BLB_UP[226] BLB_UP[227] BLEQ_DN BLEQ_UP BL_DN[224] BL_DN[225]
+ BL_DN[226] BL_DN[227] BL_UP[224] BL_UP[225] BL_UP[226] BL_UP[227] GBL[56]
+ GBLB[56] GW[56] GWB[56] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_57 BLB_DN[228] BLB_DN[229] BLB_DN[230] BLB_DN[231] BLB_UP[228]
+ BLB_UP[229] BLB_UP[230] BLB_UP[231] BLEQ_DN BLEQ_UP BL_DN[228] BL_DN[229]
+ BL_DN[230] BL_DN[231] BL_UP[228] BL_UP[229] BL_UP[230] BL_UP[231] GBL[57]
+ GBLB[57] GW[57] GWB[57] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_58 BLB_DN[232] BLB_DN[233] BLB_DN[234] BLB_DN[235] BLB_UP[232]
+ BLB_UP[233] BLB_UP[234] BLB_UP[235] BLEQ_DN BLEQ_UP BL_DN[232] BL_DN[233]
+ BL_DN[234] BL_DN[235] BL_UP[232] BL_UP[233] BL_UP[234] BL_UP[235] GBL[58]
+ GBLB[58] GW[58] GWB[58] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_59 BLB_DN[236] BLB_DN[237] BLB_DN[238] BLB_DN[239] BLB_UP[236]
+ BLB_UP[237] BLB_UP[238] BLB_UP[239] BLEQ_DN BLEQ_UP BL_DN[236] BL_DN[237]
+ BL_DN[238] BL_DN[239] BL_UP[236] BL_UP[237] BL_UP[238] BL_UP[239] GBL[59]
+ GBLB[59] GW[59] GWB[59] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_60 BLB_DN[240] BLB_DN[241] BLB_DN[242] BLB_DN[243] BLB_UP[240]
+ BLB_UP[241] BLB_UP[242] BLB_UP[243] BLEQ_DN BLEQ_UP BL_DN[240] BL_DN[241]
+ BL_DN[242] BL_DN[243] BL_UP[240] BL_UP[241] BL_UP[242] BL_UP[243] GBL[60]
+ GBLB[60] GW[60] GWB[60] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_61 BLB_DN[244] BLB_DN[245] BLB_DN[246] BLB_DN[247] BLB_UP[244]
+ BLB_UP[245] BLB_UP[246] BLB_UP[247] BLEQ_DN BLEQ_UP BL_DN[244] BL_DN[245]
+ BL_DN[246] BL_DN[247] BL_UP[244] BL_UP[245] BL_UP[246] BL_UP[247] GBL[61]
+ GBLB[61] GW[61] GWB[61] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_62 BLB_DN[248] BLB_DN[249] BLB_DN[250] BLB_DN[251] BLB_UP[248]
+ BLB_UP[249] BLB_UP[250] BLB_UP[251] BLEQ_DN BLEQ_UP BL_DN[248] BL_DN[249]
+ BL_DN[250] BL_DN[251] BL_UP[248] BL_UP[249] BL_UP[250] BL_UP[251] GBL[62]
+ GBLB[62] GW[62] GWB[62] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
XLIO_M4_63 BLB_DN[252] BLB_DN[253] BLB_DN[254] BLB_DN[255] BLB_UP[252]
+ BLB_UP[253] BLB_UP[254] BLB_UP[255] BLEQ_DN BLEQ_UP BL_DN[252] BL_DN[253]
+ BL_DN[254] BL_DN[255] BL_UP[252] BL_UP[253] BL_UP[254] BL_UP[255] GBL[63]
+ GBLB[63] GW[63] GWB[63] RE SAEB VDDHD VDDI VSSI WE YL_LIO[0] YL_LIO[1] Y_DN[0]
+ Y_DN[1] Y_DN[2] Y_DN[3] Y_DN[4] Y_DN[5] Y_DN[6] Y_DN[7] Y_UP[0] Y_UP[1]
+ Y_UP[2] Y_UP[3] Y_UP[4] Y_UP[5] Y_UP[6] Y_UP[7] S1AHSF400W40_LIO_M4
.ENDS

.SUBCKT S1AHSF400W40_BANK_F GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6]
+ GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16]
+ GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25]
+ GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34]
+ GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43]
+ GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52]
+ GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61]
+ GBL[62] GBL[63] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6]
+ GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15]
+ GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23]
+ GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31]
+ GBLB[32] GBLB[33] GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39]
+ GBLB[40] GBLB[41] GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47]
+ GBLB[48] GBLB[49] GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55]
+ GBLB[56] GBLB[57] GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3]
+ GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13]
+ GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22]
+ GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31]
+ GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40]
+ GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49]
+ GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58]
+ GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] PD_BUF PD_CVDDBUF RW_RE VDDHD WLP_SAE
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6]
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5]
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_Y[0] DEC_Y[1]
+ DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] YL[0] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] VDDI
+ VSSI WLP_SAE_TK
XLIO_MCB_F GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9]
+ GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18]
+ GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27]
+ GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36]
+ GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45]
+ GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54]
+ GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63]
+ GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8]
+ GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16]
+ GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24]
+ GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32]
+ GBLB[33] GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40]
+ GBLB[41] GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48]
+ GBLB[49] GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56]
+ GBLB[57] GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] VDDHD WL[0]
+ WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12]
+ WL[13] WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23]
+ WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34]
+ WL[35] WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45]
+ WL[46] WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56]
+ WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67]
+ WL[68] WL[69] WL[70] WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78]
+ WL[79] WL[80] WL[81] WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89]
+ WL[90] WL[91] WL[92] WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100]
+ WL[101] WL[102] WL[103] WL[104] WL[105] WL[106] WL[107] WL[108] WL[109]
+ WL[110] WL[111] WL[112] WL[113] WL[114] WL[115] WL[116] WL[117] WL[118]
+ WL[119] WL[120] WL[121] WL[122] WL[123] WL[124] WL[125] WL[126] WL[127]
+ BLEQ_DN BLEQ_UP GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9]
+ GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20]
+ GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31]
+ GW[32] GW[33] GW[34] GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42]
+ GW[43] GW[44] GW[45] GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53]
+ GW[54] GW[55] GW[56] GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] RE SAEB WE DEC_Y_DN[0]
+ DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6]
+ DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4]
+ DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] YL_LIO[0] YL_LIO[1] VDDI VSSI
+ S1AHSF400W40_LIO_MCB_F
XLCTRL_F_M4 BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4]
+ DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2]
+ DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] PD_BUF PD_CVDDBUF
+ RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] WLPY_DN[2] WLPY_DN[3]
+ WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE WLP_SAE_TK YL[0] YL_LIO[0]
+ YL_LIO[1] S1AHSF400W40_LCTRL_F_M4
XXDRV_STRAPD0 VDDHD VDDI VSSI WLPY_DN[0] WLPY_DNB[0] S1AHSF400W40_XDRV_STRAP
XXDRV_LA512_0 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[0] WL[1] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_1 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[2] WL[3] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_2 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[4] WL[5] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_3 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[6] WL[7] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_4 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[8] WL[9] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_5 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[10] WL[11] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_6 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[12] WL[13] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_7 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[14] WL[15] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_8 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[16] WL[17] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_9 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[18] WL[19] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_10 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[20] WL[21] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_11 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[22] WL[23] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_12 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[24] WL[25] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_13 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[26] WL[27] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_14 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[28] WL[29] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_15 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[30] WL[31] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_16 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[32] WL[33] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_17 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[34] WL[35] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_18 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[36] WL[37] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_19 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[38] WL[39] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_20 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[40] WL[41] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_21 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[42] WL[43] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_22 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[44] WL[45] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_23 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[46] WL[47] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_24 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[48] WL[49] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_25 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[50] WL[51] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_26 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[52] WL[53] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_27 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[54] WL[55] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_28 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[56] WL[57] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_29 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[58] WL[59] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_30 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[60] WL[61] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_31 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[62] WL[63] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_STRAPU1 VDDHD VDDI VSSI WLPY_UP[0] WLPY_UPB[0] S1AHSF400W40_XDRV_STRAP
XXDRV_LA512_32 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[64] WL[65] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_33 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[66] WL[67] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_34 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[68] WL[69] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_35 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[70] WL[71] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_36 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[72] WL[73] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_37 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[74] WL[75] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_38 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[76] WL[77] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_39 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[78] WL[79] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_40 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[80] WL[81] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_41 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[82] WL[83] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_42 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[84] WL[85] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_43 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[86] WL[87] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_44 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[88] WL[89] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_45 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[90] WL[91] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_46 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[92] WL[93] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_47 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[94] WL[95] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_48 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[96] WL[97] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_49 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[98] WL[99] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_50 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[100] WL[101] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_51 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[102] WL[103] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_52 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[104] WL[105] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_53 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[106] WL[107] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_54 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[108] WL[109] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_55 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[110] WL[111] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_56 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[112] WL[113] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_57 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[114] WL[115] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_58 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[116] WL[117] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_59 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[118] WL[119] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_60 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[120] WL[121] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_61 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[122] WL[123] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_62 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[124] WL[125] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_63 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[126] WL[127] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
.ENDS

.SUBCKT S1AHSF400W40_WL_TRK WL_TK BL_TK PD_BUF VDDHD TIEH TIEL VDDI VSSI
XTKWL_2X2_RL0 VDDI VSSI WL_TK WL_TK S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RL1 VDDI VSSI WL_TK WL_TK S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RL2 VDDI VSSI WL_TK WL_TK S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RL3 VDDI VSSI WL_TK WL_TK S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RL4 VDDI VSSI WL_TK WL_TK S1AHSF400W40_TKWL_2X2
XTKWL_2X2_ISO VDDI VSSI WL_TK WL_TK TIEL TIEL S1AHSF400W40_TKWL_2X2_ISO
XTKWL_2X2_RR0 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR1 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR2 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR3 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR4 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR5 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR6 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR7 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR8 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR9 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR10 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR11 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR12 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR13 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR14 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR15 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR16 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR17 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR18 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR19 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR20 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR21 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR22 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR23 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR24 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR25 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR26 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR27 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR28 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR29 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR30 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR31 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR32 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR33 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR34 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR35 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR36 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR37 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR38 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR39 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR40 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR41 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR42 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR43 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR44 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR45 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR46 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR47 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR48 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR49 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR50 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR51 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR52 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR53 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR54 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR55 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR56 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR57 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_RR58 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKBL_TRKPRE PD_BUF BL_TK WL_TK VDDHD VDDI VSSI TIEH TIEL
+ S1AHSF400W40_TKBL_TRKPRE
XTKWL_2X2_L0 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L1 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L2 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L3 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L4 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L5 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L6 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L7 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L8 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L9 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L10 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L11 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L12 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L13 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L14 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L15 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L16 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L17 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L18 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L19 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L20 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L21 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L22 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L23 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L24 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L25 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L26 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L27 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L28 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L29 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L30 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L31 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L32 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L33 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L34 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L35 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L36 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L37 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L38 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L39 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L40 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L41 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L42 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L43 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L44 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L45 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L46 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L47 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L48 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L49 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L50 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L51 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L52 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L53 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L54 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L55 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L56 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L57 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L58 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L59 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L60 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L61 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L62 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
XTKWL_2X2_L63 VDDI VSSI TIEL TIEL S1AHSF400W40_TKWL_2X2
.ENDS

.SUBCKT S1AHSF400W40_TRACKING WL_TK PD_BUF BL_TK VDDHD WL[0] WL[1] WL[2] WL[3]
+ WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15]
+ WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26]
+ WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37]
+ WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48]
+ WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59]
+ WL[60] WL[61] WL[62] WL[63] VDDI VSSI
XWL_TRK WL_TK BL_TK PD_BUF VDDHD TIEH TIEL VDDI VSSI S1AHSF400W40_WL_TRK
X0TRKNORX2_0 BL_TK VDDI VSSI WL[0] WL[1] WL_TK FLOAT1[0] NET[0] FLOAT3 FLOAT4[0]
+ TIEH S1AHSF400W40_TRKNORX2
X1TRKNORX2_1 BL_TK VDDI VSSI WL[2] WL[3] WL_TK FLOAT1[1] NET[1] NET[0] FLOAT4[1]
+ TIEH S1AHSF400W40_TRKNORX2
X2TRKNORX2_2 BL_TK VDDI VSSI WL[4] WL[5] WL_TK FLOAT1[2] NET[2] NET[1] FLOAT4[2]
+ TIEH S1AHSF400W40_TRKNORX2
X3TRKNORX2_3 BL_TK VDDI VSSI WL[6] WL[7] WL_TK FLOAT1[3] NET[3] NET[2] FLOAT4[3]
+ TIEH S1AHSF400W40_TRKNORX2
X2TRKNORX2_4 BL_TK VDDI VSSI WL[8] WL[9] WL_TK FLOAT1[4] NET[4] NET[3] FLOAT4[4]
+ TIEH S1AHSF400W40_TRKNORX2
X3TRKNORX2_5 BL_TK VDDI VSSI WL[10] WL[11] WL_TK FLOAT1[5] NET[5] NET[4]
+ FLOAT4[5] TIEH S1AHSF400W40_TRKNORX2
X2TRKNORX2_6 BL_TK VDDI VSSI WL[12] WL[13] WL_TK FLOAT1[6] NET[6] NET[5]
+ FLOAT4[6] TIEH S1AHSF400W40_TRKNORX2
X3TRKNORX2_7 BL_TK VDDI VSSI WL[14] WL[15] WL_TK FLOAT1[7] NET[7] NET[6]
+ FLOAT4[7] TIEH S1AHSF400W40_TRKNORX2
X2TRKNORX2_8 BL_TK VDDI VSSI WL[16] WL[17] WL_TK FLOAT1[8] NET[8] NET[7]
+ FLOAT4[8] TIEH S1AHSF400W40_TRKNORX2
X3TRKNORX2_9 BL_TK VDDI VSSI WL[18] WL[19] WL_TK FLOAT1[9] NET[9] NET[8]
+ FLOAT4[9] TIEH S1AHSF400W40_TRKNORX2
X2TRKNORX2_10 BL_TK VDDI VSSI WL[20] WL[21] WL_TK FLOAT1[10] NET[10] NET[9]
+ FLOAT4[10] TIEH S1AHSF400W40_TRKNORX2
X3TRKNORX2_11 BL_TK VDDI VSSI WL[22] WL[23] WL_TK FLOAT1[11] NET[11] NET[10]
+ FLOAT4[11] TIEH S1AHSF400W40_TRKNORX2
X2TRKNORX2_12 BL_TK VDDI VSSI WL[24] WL[25] WL_TK FLOAT1[12] NET[12] NET[11]
+ FLOAT4[12] TIEH S1AHSF400W40_TRKNORX2
X3TRKNORX2_13 BL_TK VDDI VSSI WL[26] WL[27] WL_TK FLOAT1[13] NET[13] NET[12]
+ FLOAT4[13] TIEH S1AHSF400W40_TRKNORX2
X2TRKNORX2_14 BL_TK VDDI VSSI WL[28] WL[29] WL_TK FLOAT1[14] NET[14] NET[13]
+ FLOAT4[14] TIEH S1AHSF400W40_TRKNORX2
X3TRKNORX2_15 BL_TK VDDI VSSI WL[30] WL[31] WL_TK FLOAT1[15] NET[15] NET[14]
+ FLOAT4[15] TIEH S1AHSF400W40_TRKNORX2
X2TRKNORX2_16 BL_TK VDDI VSSI WL[32] WL[33] WL_TK FLOAT1[16] NET[16] NET[15]
+ FLOAT4[16] TIEH S1AHSF400W40_TRKNORX2
X3TRKNORX2_17 BL_TK VDDI VSSI WL[34] WL[35] WL_TK FLOAT1[17] NET[17] NET[16]
+ FLOAT4[17] TIEH S1AHSF400W40_TRKNORX2
X2TRKNORX2_18 BL_TK VDDI VSSI WL[36] WL[37] WL_TK FLOAT1[18] NET[18] NET[17]
+ FLOAT4[18] TIEH S1AHSF400W40_TRKNORX2
X3TRKNORX2_19 BL_TK VDDI VSSI WL[38] WL[39] WL_TK FLOAT1[19] NET[19] NET[18]
+ FLOAT4[19] TIEH S1AHSF400W40_TRKNORX2
X2TRKNORX2_20 BL_TK VDDI VSSI WL[40] WL[41] WL_TK FLOAT1[20] NET[20] NET[19]
+ FLOAT4[20] TIEH S1AHSF400W40_TRKNORX2
X3TRKNORX2_21 BL_TK VDDI VSSI WL[42] WL[43] WL_TK FLOAT1[21] NET[21] NET[20]
+ FLOAT4[21] TIEH S1AHSF400W40_TRKNORX2
X2TRKNORX2_22 BL_TK VDDI VSSI WL[44] WL[45] WL_TK FLOAT1[22] NET[22] NET[21]
+ FLOAT4[22] TIEH S1AHSF400W40_TRKNORX2
X3TRKNORX2_23 BL_TK VDDI VSSI WL[46] WL[47] WL_TK FLOAT1[23] NET[23] NET[22]
+ FLOAT4[23] TIEH S1AHSF400W40_TRKNORX2
X2TRKNORX2_24 BL_TK VDDI VSSI WL[48] WL[49] WL_TK FLOAT1[24] NET[24] NET[23]
+ FLOAT4[24] TIEH S1AHSF400W40_TRKNORX2
X3TRKNORX2_25 BL_TK VDDI VSSI WL[50] WL[51] WL_TK FLOAT1[25] NET[25] NET[24]
+ FLOAT4[25] TIEH S1AHSF400W40_TRKNORX2
X2TRKNORX2_26 BL_TK VDDI VSSI WL[52] WL[53] WL_TK FLOAT1[26] NET[26] NET[25]
+ FLOAT4[26] TIEH S1AHSF400W40_TRKNORX2
X3TRKNORX2_27 BL_TK VDDI VSSI WL[54] WL[55] WL_TK FLOAT1[27] NET[27] NET[26]
+ FLOAT4[27] TIEH S1AHSF400W40_TRKNORX2
X2TRKNORX2_28 BL_TK VDDI VSSI WL[56] WL[57] WL_TK FLOAT1[28] NET[28] NET[27]
+ FLOAT4[28] TIEH S1AHSF400W40_TRKNORX2
X3TRKNORX2_29 BL_TK VDDI VSSI WL[58] WL[59] WL_TK FLOAT1[29] NET[29] NET[28]
+ FLOAT4[29] TIEH S1AHSF400W40_TRKNORX2
X2TRKNORX2_30 BL_TK VDDI VSSI WL[60] WL[61] WL_TK FLOAT1[30] NET[30] NET[29]
+ FLOAT4[30] TIEH S1AHSF400W40_TRKNORX2
X3TRKNORX2_31 BL_TK VDDI VSSI WL[62] WL[63] WL_TK FLOAT1[31] NET[31] NET[30]
+ FLOAT4[31] TIEH S1AHSF400W40_TRKNORX2
.ENDS

.SUBCKT S1AHSF400W40_BANK_0_F GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6]
+ GBL[7] GBL[8] GBL[9] GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16]
+ GBL[17] GBL[18] GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25]
+ GBL[26] GBL[27] GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34]
+ GBL[35] GBL[36] GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43]
+ GBL[44] GBL[45] GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52]
+ GBL[53] GBL[54] GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61]
+ GBL[62] GBL[63] GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6]
+ GBLB[7] GBLB[8] GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15]
+ GBLB[16] GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23]
+ GBLB[24] GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31]
+ GBLB[32] GBLB[33] GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39]
+ GBLB[40] GBLB[41] GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47]
+ GBLB[48] GBLB[49] GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55]
+ GBLB[56] GBLB[57] GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0]
+ GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12]
+ GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23]
+ GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34]
+ GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45]
+ GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56]
+ GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3]
+ GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13]
+ GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22]
+ GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31]
+ GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40]
+ GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49]
+ GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58]
+ GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] PD_BUF PD_CVDDBUF RW_RE VDDHD WLP_SAE
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6]
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5]
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_Y[0] DEC_Y[1]
+ DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] YL[0] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] BL_TK
+ WL_TK VDDI VSSI WLP_SAE_TK
XTRACKING WL_TK PD_BUF BL_TK VDDHD WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6]
+ WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17]
+ WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28]
+ WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39]
+ WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50]
+ WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61]
+ WL[62] WL[63] VDDI VSSI S1AHSF400W40_TRACKING
XLIO_MCB_F GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9]
+ GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18]
+ GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27]
+ GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36]
+ GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45]
+ GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54]
+ GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63]
+ GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8]
+ GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16]
+ GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24]
+ GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32]
+ GBLB[33] GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40]
+ GBLB[41] GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48]
+ GBLB[49] GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56]
+ GBLB[57] GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] VDDHD WL[0]
+ WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12]
+ WL[13] WL[14] WL[15] WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23]
+ WL[24] WL[25] WL[26] WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34]
+ WL[35] WL[36] WL[37] WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45]
+ WL[46] WL[47] WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56]
+ WL[57] WL[58] WL[59] WL[60] WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67]
+ WL[68] WL[69] WL[70] WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78]
+ WL[79] WL[80] WL[81] WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89]
+ WL[90] WL[91] WL[92] WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100]
+ WL[101] WL[102] WL[103] WL[104] WL[105] WL[106] WL[107] WL[108] WL[109]
+ WL[110] WL[111] WL[112] WL[113] WL[114] WL[115] WL[116] WL[117] WL[118]
+ WL[119] WL[120] WL[121] WL[122] WL[123] WL[124] WL[125] WL[126] WL[127]
+ BLEQ_DN BLEQ_UP GW[0] GW[1] GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9]
+ GW[10] GW[11] GW[12] GW[13] GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20]
+ GW[21] GW[22] GW[23] GW[24] GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31]
+ GW[32] GW[33] GW[34] GW[35] GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42]
+ GW[43] GW[44] GW[45] GW[46] GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53]
+ GW[54] GW[55] GW[56] GW[57] GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GWB[0]
+ GWB[1] GWB[2] GWB[3] GWB[4] GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11]
+ GWB[12] GWB[13] GWB[14] GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20]
+ GWB[21] GWB[22] GWB[23] GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29]
+ GWB[30] GWB[31] GWB[32] GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38]
+ GWB[39] GWB[40] GWB[41] GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47]
+ GWB[48] GWB[49] GWB[50] GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56]
+ GWB[57] GWB[58] GWB[59] GWB[60] GWB[61] GWB[62] GWB[63] RE SAEB WE DEC_Y_DN[0]
+ DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4] DEC_Y_DN[5] DEC_Y_DN[6]
+ DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2] DEC_Y_UP[3] DEC_Y_UP[4]
+ DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] YL_LIO[0] YL_LIO[1] VDDI VSSI
+ S1AHSF400W40_LIO_MCB_F
XLCTRL_F_M4 BLEQ_DN BLEQ_UP DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4]
+ DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2]
+ DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5]
+ DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5]
+ DEC_Y[6] DEC_Y[7] DEC_Y_DN[0] DEC_Y_DN[1] DEC_Y_DN[2] DEC_Y_DN[3] DEC_Y_DN[4]
+ DEC_Y_DN[5] DEC_Y_DN[6] DEC_Y_DN[7] DEC_Y_UP[0] DEC_Y_UP[1] DEC_Y_UP[2]
+ DEC_Y_UP[3] DEC_Y_UP[4] DEC_Y_UP[5] DEC_Y_UP[6] DEC_Y_UP[7] PD_BUF PD_CVDDBUF
+ RE RW_RE SAEB VDDHD VDDI VSSI WE WLPY_DN[0] WLPY_DN[1] WLPY_DN[2] WLPY_DN[3]
+ WLPY_UP[0] WLPY_UP[1] WLPY_UP[2] WLPY_UP[3] WLP_SAE WLP_SAE_TK YL[0] YL_LIO[0]
+ YL_LIO[1] S1AHSF400W40_LCTRL_F_M4
XXDRV_STRAPD0 VDDHD VDDI VSSI WLPY_DN[0] WLPY_DNB[0] S1AHSF400W40_XDRV_STRAP
XXDRV_LA512_0 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[0] WL[1] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_1 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[2] WL[3] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_2 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[4] WL[5] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_3 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[6] WL[7] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_4 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[8] WL[9] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_5 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[10] WL[11] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_6 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[12] WL[13] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_7 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[14] WL[15] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_8 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[16] WL[17] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_9 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[18] WL[19] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_10 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[20] WL[21] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_11 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[22] WL[23] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_12 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[24] WL[25] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_13 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[26] WL[27] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_14 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[28] WL[29] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_15 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[30] WL[31] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_16 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[32] WL[33] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_17 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[34] WL[35] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_18 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[36] WL[37] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_19 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[38] WL[39] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_20 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[40] WL[41] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_21 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[42] WL[43] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_22 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[44] WL[45] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_23 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[46] WL[47] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_24 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[48] WL[49] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_25 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[50] WL[51] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_26 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[52] WL[53] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_27 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[54] WL[55] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_28 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[56] WL[57] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_29 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[58] WL[59] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_30 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[60] WL[61] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_31 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[62] WL[63] WLPY_DN[0]
+ WLPY_DNB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_STRAPU1 VDDHD VDDI VSSI WLPY_UP[0] WLPY_UPB[0] S1AHSF400W40_XDRV_STRAP
XXDRV_LA512_32 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[64] WL[65] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_33 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[66] WL[67] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_34 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[68] WL[69] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_35 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[70] WL[71] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_36 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[72] WL[73] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_37 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[74] WL[75] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_38 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[76] WL[77] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_39 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[1] DEC_X1[0] DEC_X1[2] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[78] WL[79] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_40 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[80] WL[81] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_41 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[82] WL[83] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_42 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[84] WL[85] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_43 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[2] DEC_X1[0] DEC_X1[1] DEC_X1[3] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[86] WL[87] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_44 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[88] WL[89] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_45 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[90] WL[91] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_46 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[92] WL[93] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_47 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[3] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[4]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[94] WL[95] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_48 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[96] WL[97] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_49 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[98] WL[99] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_50 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[100] WL[101] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_51 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[4] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[5] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[102] WL[103] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_52 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[104] WL[105] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_53 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[106] WL[107] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_54 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[108] WL[109] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_55 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[5] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[110] WL[111] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_56 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[112] WL[113] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_57 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[114] WL[115] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_58 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[116] WL[117] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_59 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[6] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[118] WL[119] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_60 DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[120] WL[121] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_61 DEC_X0[2] DEC_X0[3] DEC_X0[0] DEC_X0[1] DEC_X0[4] DEC_X0[5]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[122] WL[123] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_62 DEC_X0[4] DEC_X0[5] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[6] DEC_X0[7] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[124] WL[125] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
XXDRV_LA512_63 DEC_X0[6] DEC_X0[7] DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3]
+ DEC_X0[4] DEC_X0[5] DEC_X1[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3]
+ DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3]
+ DEC_X3[0] DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6]
+ DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6]
+ DEC_Y[7] PD_BUF PD_CVDDBUF RW_RE VDDHD VDDI VSSI WL[126] WL[127] WLPY_UP[0]
+ WLPY_UPB[0] WLP_SAE WLP_SAE_TK YL[0] S1AHSF400W40_XDRV_LA512
.ENDS

.SUBCKT TS1N65LPHSA1024X64M4F Q[63] Q[62] Q[61] Q[60] Q[59] Q[58] Q[57] Q[56]
+ Q[55] Q[54] Q[53] Q[52] Q[51] Q[50] Q[49] Q[48] Q[47] Q[46] Q[45] Q[44] Q[43]
+ Q[42] Q[41] Q[40] Q[39] Q[38] Q[37] Q[36] Q[35] Q[34] Q[33] Q[32] Q[31] Q[30]
+ Q[29] Q[28] Q[27] Q[26] Q[25] Q[24] Q[23] Q[22] Q[21] Q[20] Q[19] Q[18] Q[17]
+ Q[16] Q[15] Q[14] Q[13] Q[12] Q[11] Q[10] Q[9] Q[8] Q[7] Q[6] Q[5] Q[4] Q[3]
+ Q[2] Q[1] Q[0] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] BWEB[63]
+ BWEB[62] BWEB[61] BWEB[60] BWEB[59] BWEB[58] BWEB[57] BWEB[56] BWEB[55]
+ BWEB[54] BWEB[53] BWEB[52] BWEB[51] BWEB[50] BWEB[49] BWEB[48] BWEB[47]
+ BWEB[46] BWEB[45] BWEB[44] BWEB[43] BWEB[42] BWEB[41] BWEB[40] BWEB[39]
+ BWEB[38] BWEB[37] BWEB[36] BWEB[35] BWEB[34] BWEB[33] BWEB[32] BWEB[31]
+ BWEB[30] BWEB[29] BWEB[28] BWEB[27] BWEB[26] BWEB[25] BWEB[24] BWEB[23]
+ BWEB[22] BWEB[21] BWEB[20] BWEB[19] BWEB[18] BWEB[17] BWEB[16] BWEB[15]
+ BWEB[14] BWEB[13] BWEB[12] BWEB[11] BWEB[10] BWEB[9] BWEB[8] BWEB[7] BWEB[6]
+ BWEB[5] BWEB[4] BWEB[3] BWEB[2] BWEB[1] BWEB[0] CEB CLK D[63] D[62] D[61]
+ D[60] D[59] D[58] D[57] D[56] D[55] D[54] D[53] D[52] D[51] D[50] D[49] D[48]
+ D[47] D[46] D[45] D[44] D[43] D[42] D[41] D[40] D[39] D[38] D[37] D[36] D[35]
+ D[34] D[33] D[32] D[31] D[30] D[29] D[28] D[27] D[26] D[25] D[24] D[23] D[22]
+ D[21] D[20] D[19] D[18] D[17] D[16] D[15] D[14] D[13] D[12] D[11] D[10] D[9]
+ D[8] D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] RTSEL[1] RTSEL[0] WTSEL[2]
+ WTSEL[1] WTSEL[0] WEB VDD VSS
XBANK_S_0 GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9]
+ GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18]
+ GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27]
+ GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36]
+ GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45]
+ GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54]
+ GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63]
+ GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8]
+ GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16]
+ GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24]
+ GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32]
+ GBLB[33] GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40]
+ GBLB[41] GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48]
+ GBLB[49] GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56]
+ GBLB[57] GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1]
+ GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13]
+ GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24]
+ GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35]
+ GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46]
+ GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57]
+ GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4]
+ GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14]
+ GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23]
+ GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32]
+ GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41]
+ GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50]
+ GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59]
+ GWB[60] GWB[61] GWB[62] GWB[63] PD_BUF PD_CVDDBUF RW_RE VDDHD WLP_SAE
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6]
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5]
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_Y[0] DEC_Y[1]
+ DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] YL[0] DEC_X3[0]
+ DEC_X3[1] DEC_X3[2] DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] TRKBL
+ BLTRKWLDRV VDD VSS WLP_SAE_TK S1AHSF400W40_BANK_0_F
XBANK_S_1 GBL[0] GBL[1] GBL[2] GBL[3] GBL[4] GBL[5] GBL[6] GBL[7] GBL[8] GBL[9]
+ GBL[10] GBL[11] GBL[12] GBL[13] GBL[14] GBL[15] GBL[16] GBL[17] GBL[18]
+ GBL[19] GBL[20] GBL[21] GBL[22] GBL[23] GBL[24] GBL[25] GBL[26] GBL[27]
+ GBL[28] GBL[29] GBL[30] GBL[31] GBL[32] GBL[33] GBL[34] GBL[35] GBL[36]
+ GBL[37] GBL[38] GBL[39] GBL[40] GBL[41] GBL[42] GBL[43] GBL[44] GBL[45]
+ GBL[46] GBL[47] GBL[48] GBL[49] GBL[50] GBL[51] GBL[52] GBL[53] GBL[54]
+ GBL[55] GBL[56] GBL[57] GBL[58] GBL[59] GBL[60] GBL[61] GBL[62] GBL[63]
+ GBLB[0] GBLB[1] GBLB[2] GBLB[3] GBLB[4] GBLB[5] GBLB[6] GBLB[7] GBLB[8]
+ GBLB[9] GBLB[10] GBLB[11] GBLB[12] GBLB[13] GBLB[14] GBLB[15] GBLB[16]
+ GBLB[17] GBLB[18] GBLB[19] GBLB[20] GBLB[21] GBLB[22] GBLB[23] GBLB[24]
+ GBLB[25] GBLB[26] GBLB[27] GBLB[28] GBLB[29] GBLB[30] GBLB[31] GBLB[32]
+ GBLB[33] GBLB[34] GBLB[35] GBLB[36] GBLB[37] GBLB[38] GBLB[39] GBLB[40]
+ GBLB[41] GBLB[42] GBLB[43] GBLB[44] GBLB[45] GBLB[46] GBLB[47] GBLB[48]
+ GBLB[49] GBLB[50] GBLB[51] GBLB[52] GBLB[53] GBLB[54] GBLB[55] GBLB[56]
+ GBLB[57] GBLB[58] GBLB[59] GBLB[60] GBLB[61] GBLB[62] GBLB[63] GW[0] GW[1]
+ GW[2] GW[3] GW[4] GW[5] GW[6] GW[7] GW[8] GW[9] GW[10] GW[11] GW[12] GW[13]
+ GW[14] GW[15] GW[16] GW[17] GW[18] GW[19] GW[20] GW[21] GW[22] GW[23] GW[24]
+ GW[25] GW[26] GW[27] GW[28] GW[29] GW[30] GW[31] GW[32] GW[33] GW[34] GW[35]
+ GW[36] GW[37] GW[38] GW[39] GW[40] GW[41] GW[42] GW[43] GW[44] GW[45] GW[46]
+ GW[47] GW[48] GW[49] GW[50] GW[51] GW[52] GW[53] GW[54] GW[55] GW[56] GW[57]
+ GW[58] GW[59] GW[60] GW[61] GW[62] GW[63] GWB[0] GWB[1] GWB[2] GWB[3] GWB[4]
+ GWB[5] GWB[6] GWB[7] GWB[8] GWB[9] GWB[10] GWB[11] GWB[12] GWB[13] GWB[14]
+ GWB[15] GWB[16] GWB[17] GWB[18] GWB[19] GWB[20] GWB[21] GWB[22] GWB[23]
+ GWB[24] GWB[25] GWB[26] GWB[27] GWB[28] GWB[29] GWB[30] GWB[31] GWB[32]
+ GWB[33] GWB[34] GWB[35] GWB[36] GWB[37] GWB[38] GWB[39] GWB[40] GWB[41]
+ GWB[42] GWB[43] GWB[44] GWB[45] GWB[46] GWB[47] GWB[48] GWB[49] GWB[50]
+ GWB[51] GWB[52] GWB[53] GWB[54] GWB[55] GWB[56] GWB[57] GWB[58] GWB[59]
+ GWB[60] GWB[61] GWB[62] GWB[63] PD_BUF PD_CVDDBUF RW_RE VDDHD WLP_SAE
+ DEC_X0[0] DEC_X0[1] DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6]
+ DEC_X0[7] DEC_X1[0] DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5]
+ DEC_X1[6] DEC_X1[7] DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_Y[0] DEC_Y[1]
+ DEC_Y[2] DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] YL[0] DEC_X3[2]
+ DEC_X3[3] DEC_X3[0] DEC_X3[1] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] VDD VSS
+ WLP_SAE_TK S1AHSF400W40_BANK_F
XIO_M4_0 AWT2 BIST2IO BWEB[0] VLO CKD D[0] VLO GBL[0] GBLB[0] GW[0] GWB[0]
+ PD_BUF Q[0] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_1 AWT2 BIST2IO BWEB[1] VLO CKD D[1] VLO GBL[1] GBLB[1] GW[1] GWB[1]
+ PD_BUF Q[1] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_2 AWT2 BIST2IO BWEB[2] VLO CKD D[2] VLO GBL[2] GBLB[2] GW[2] GWB[2]
+ PD_BUF Q[2] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_3 AWT2 BIST2IO BWEB[3] VLO CKD D[3] VLO GBL[3] GBLB[3] GW[3] GWB[3]
+ PD_BUF Q[3] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_4 AWT2 BIST2IO BWEB[4] VLO CKD D[4] VLO GBL[4] GBLB[4] GW[4] GWB[4]
+ PD_BUF Q[4] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_5 AWT2 BIST2IO BWEB[5] VLO CKD D[5] VLO GBL[5] GBLB[5] GW[5] GWB[5]
+ PD_BUF Q[5] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_6 AWT2 BIST2IO BWEB[6] VLO CKD D[6] VLO GBL[6] GBLB[6] GW[6] GWB[6]
+ PD_BUF Q[6] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_7 AWT2 BIST2IO BWEB[7] VLO CKD D[7] VLO GBL[7] GBLB[7] GW[7] GWB[7]
+ PD_BUF Q[7] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_8 AWT2 BIST2IO BWEB[8] VLO CKD D[8] VLO GBL[8] GBLB[8] GW[8] GWB[8]
+ PD_BUF Q[8] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_9 AWT2 BIST2IO BWEB[9] VLO CKD D[9] VLO GBL[9] GBLB[9] GW[9] GWB[9]
+ PD_BUF Q[9] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_10 AWT2 BIST2IO BWEB[10] VLO CKD D[10] VLO GBL[10] GBLB[10] GW[10]
+ GWB[10] PD_BUF Q[10] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_11 AWT2 BIST2IO BWEB[11] VLO CKD D[11] VLO GBL[11] GBLB[11] GW[11]
+ GWB[11] PD_BUF Q[11] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_12 AWT2 BIST2IO BWEB[12] VLO CKD D[12] VLO GBL[12] GBLB[12] GW[12]
+ GWB[12] PD_BUF Q[12] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_13 AWT2 BIST2IO BWEB[13] VLO CKD D[13] VLO GBL[13] GBLB[13] GW[13]
+ GWB[13] PD_BUF Q[13] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_14 AWT2 BIST2IO BWEB[14] VLO CKD D[14] VLO GBL[14] GBLB[14] GW[14]
+ GWB[14] PD_BUF Q[14] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_15 AWT2 BIST2IO BWEB[15] VLO CKD D[15] VLO GBL[15] GBLB[15] GW[15]
+ GWB[15] PD_BUF Q[15] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_16 AWT2 BIST2IO BWEB[16] VLO CKD D[16] VLO GBL[16] GBLB[16] GW[16]
+ GWB[16] PD_BUF Q[16] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_17 AWT2 BIST2IO BWEB[17] VLO CKD D[17] VLO GBL[17] GBLB[17] GW[17]
+ GWB[17] PD_BUF Q[17] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_18 AWT2 BIST2IO BWEB[18] VLO CKD D[18] VLO GBL[18] GBLB[18] GW[18]
+ GWB[18] PD_BUF Q[18] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_19 AWT2 BIST2IO BWEB[19] VLO CKD D[19] VLO GBL[19] GBLB[19] GW[19]
+ GWB[19] PD_BUF Q[19] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_20 AWT2 BIST2IO BWEB[20] VLO CKD D[20] VLO GBL[20] GBLB[20] GW[20]
+ GWB[20] PD_BUF Q[20] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_21 AWT2 BIST2IO BWEB[21] VLO CKD D[21] VLO GBL[21] GBLB[21] GW[21]
+ GWB[21] PD_BUF Q[21] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_22 AWT2 BIST2IO BWEB[22] VLO CKD D[22] VLO GBL[22] GBLB[22] GW[22]
+ GWB[22] PD_BUF Q[22] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_23 AWT2 BIST2IO BWEB[23] VLO CKD D[23] VLO GBL[23] GBLB[23] GW[23]
+ GWB[23] PD_BUF Q[23] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_24 AWT2 BIST2IO BWEB[24] VLO CKD D[24] VLO GBL[24] GBLB[24] GW[24]
+ GWB[24] PD_BUF Q[24] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_25 AWT2 BIST2IO BWEB[25] VLO CKD D[25] VLO GBL[25] GBLB[25] GW[25]
+ GWB[25] PD_BUF Q[25] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_26 AWT2 BIST2IO BWEB[26] VLO CKD D[26] VLO GBL[26] GBLB[26] GW[26]
+ GWB[26] PD_BUF Q[26] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_27 AWT2 BIST2IO BWEB[27] VLO CKD D[27] VLO GBL[27] GBLB[27] GW[27]
+ GWB[27] PD_BUF Q[27] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_28 AWT2 BIST2IO BWEB[28] VLO CKD D[28] VLO GBL[28] GBLB[28] GW[28]
+ GWB[28] PD_BUF Q[28] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_29 AWT2 BIST2IO BWEB[29] VLO CKD D[29] VLO GBL[29] GBLB[29] GW[29]
+ GWB[29] PD_BUF Q[29] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_30 AWT2 BIST2IO BWEB[30] VLO CKD D[30] VLO GBL[30] GBLB[30] GW[30]
+ GWB[30] PD_BUF Q[30] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_31 AWT2 BIST2IO BWEB[31] VLO CKD D[31] VLO GBL[31] GBLB[31] GW[31]
+ GWB[31] PD_BUF Q[31] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_32 AWT2 BIST2IO BWEB[32] VLO CKD D[32] VLO GBL[32] GBLB[32] GW[32]
+ GWB[32] PD_BUF Q[32] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_33 AWT2 BIST2IO BWEB[33] VLO CKD D[33] VLO GBL[33] GBLB[33] GW[33]
+ GWB[33] PD_BUF Q[33] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_34 AWT2 BIST2IO BWEB[34] VLO CKD D[34] VLO GBL[34] GBLB[34] GW[34]
+ GWB[34] PD_BUF Q[34] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_35 AWT2 BIST2IO BWEB[35] VLO CKD D[35] VLO GBL[35] GBLB[35] GW[35]
+ GWB[35] PD_BUF Q[35] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_36 AWT2 BIST2IO BWEB[36] VLO CKD D[36] VLO GBL[36] GBLB[36] GW[36]
+ GWB[36] PD_BUF Q[36] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_37 AWT2 BIST2IO BWEB[37] VLO CKD D[37] VLO GBL[37] GBLB[37] GW[37]
+ GWB[37] PD_BUF Q[37] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_38 AWT2 BIST2IO BWEB[38] VLO CKD D[38] VLO GBL[38] GBLB[38] GW[38]
+ GWB[38] PD_BUF Q[38] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_39 AWT2 BIST2IO BWEB[39] VLO CKD D[39] VLO GBL[39] GBLB[39] GW[39]
+ GWB[39] PD_BUF Q[39] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_40 AWT2 BIST2IO BWEB[40] VLO CKD D[40] VLO GBL[40] GBLB[40] GW[40]
+ GWB[40] PD_BUF Q[40] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_41 AWT2 BIST2IO BWEB[41] VLO CKD D[41] VLO GBL[41] GBLB[41] GW[41]
+ GWB[41] PD_BUF Q[41] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_42 AWT2 BIST2IO BWEB[42] VLO CKD D[42] VLO GBL[42] GBLB[42] GW[42]
+ GWB[42] PD_BUF Q[42] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_43 AWT2 BIST2IO BWEB[43] VLO CKD D[43] VLO GBL[43] GBLB[43] GW[43]
+ GWB[43] PD_BUF Q[43] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_44 AWT2 BIST2IO BWEB[44] VLO CKD D[44] VLO GBL[44] GBLB[44] GW[44]
+ GWB[44] PD_BUF Q[44] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_45 AWT2 BIST2IO BWEB[45] VLO CKD D[45] VLO GBL[45] GBLB[45] GW[45]
+ GWB[45] PD_BUF Q[45] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_46 AWT2 BIST2IO BWEB[46] VLO CKD D[46] VLO GBL[46] GBLB[46] GW[46]
+ GWB[46] PD_BUF Q[46] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_47 AWT2 BIST2IO BWEB[47] VLO CKD D[47] VLO GBL[47] GBLB[47] GW[47]
+ GWB[47] PD_BUF Q[47] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_48 AWT2 BIST2IO BWEB[48] VLO CKD D[48] VLO GBL[48] GBLB[48] GW[48]
+ GWB[48] PD_BUF Q[48] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_49 AWT2 BIST2IO BWEB[49] VLO CKD D[49] VLO GBL[49] GBLB[49] GW[49]
+ GWB[49] PD_BUF Q[49] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_50 AWT2 BIST2IO BWEB[50] VLO CKD D[50] VLO GBL[50] GBLB[50] GW[50]
+ GWB[50] PD_BUF Q[50] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_51 AWT2 BIST2IO BWEB[51] VLO CKD D[51] VLO GBL[51] GBLB[51] GW[51]
+ GWB[51] PD_BUF Q[51] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_52 AWT2 BIST2IO BWEB[52] VLO CKD D[52] VLO GBL[52] GBLB[52] GW[52]
+ GWB[52] PD_BUF Q[52] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_53 AWT2 BIST2IO BWEB[53] VLO CKD D[53] VLO GBL[53] GBLB[53] GW[53]
+ GWB[53] PD_BUF Q[53] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_54 AWT2 BIST2IO BWEB[54] VLO CKD D[54] VLO GBL[54] GBLB[54] GW[54]
+ GWB[54] PD_BUF Q[54] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_55 AWT2 BIST2IO BWEB[55] VLO CKD D[55] VLO GBL[55] GBLB[55] GW[55]
+ GWB[55] PD_BUF Q[55] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_56 AWT2 BIST2IO BWEB[56] VLO CKD D[56] VLO GBL[56] GBLB[56] GW[56]
+ GWB[56] PD_BUF Q[56] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_57 AWT2 BIST2IO BWEB[57] VLO CKD D[57] VLO GBL[57] GBLB[57] GW[57]
+ GWB[57] PD_BUF Q[57] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_58 AWT2 BIST2IO BWEB[58] VLO CKD D[58] VLO GBL[58] GBLB[58] GW[58]
+ GWB[58] PD_BUF Q[58] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_59 AWT2 BIST2IO BWEB[59] VLO CKD D[59] VLO GBL[59] GBLB[59] GW[59]
+ GWB[59] PD_BUF Q[59] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_60 AWT2 BIST2IO BWEB[60] VLO CKD D[60] VLO GBL[60] GBLB[60] GW[60]
+ GWB[60] PD_BUF Q[60] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_61 AWT2 BIST2IO BWEB[61] VLO CKD D[61] VLO GBL[61] GBLB[61] GW[61]
+ GWB[61] PD_BUF Q[61] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_62 AWT2 BIST2IO BWEB[62] VLO CKD D[62] VLO GBL[62] GBLB[62] GW[62]
+ GWB[62] PD_BUF Q[62] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XIO_M4_63 AWT2 BIST2IO BWEB[63] VLO CKD D[63] VLO GBL[63] GBLB[63] GW[63]
+ GWB[63] PD_BUF Q[63] VDDHD VDD VSS WLP_SAEB S1AHSF400W40_IO_M4
XCNT_CORE_M4 VLO AWT2 VLO BIST2IO BLTRKWLDRV CEB VLO CKD CLK DEC_X0[0] DEC_X0[1]
+ DEC_X0[2] DEC_X0[3] DEC_X0[4] DEC_X0[5] DEC_X0[6] DEC_X0[7] DEC_X1[0]
+ DEC_X1[1] DEC_X1[2] DEC_X1[3] DEC_X1[4] DEC_X1[5] DEC_X1[6] DEC_X1[7]
+ DEC_X2[0] DEC_X2[1] DEC_X2[2] DEC_X2[3] DEC_X3[0] DEC_X3[1] DEC_X3[2]
+ DEC_X3[3] DEC_X3[4] DEC_X3[5] DEC_X3[6] DEC_X3[7] DEC_Y[0] DEC_Y[1] DEC_Y[2]
+ DEC_Y[3] DEC_Y[4] DEC_Y[5] DEC_Y[6] DEC_Y[7] VLO PD_BUF PD_CVDDBUF PTSEL VLO
+ VLO RTSEL[0] RTSEL[1] RW_RE TK VLO TRKBL VDDHD VDD VHI VLO VSS WEB VLO WLP_SAE
+ WLP_SAEB WLP_SAE_TK WTSEL[0] WTSEL[1] WTSEL[2] A[2] A[3] A[4] A[5] A[6] A[7]
+ VLO VLO A[8] A[9] VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO VLO A[0] A[1]
+ VLO VLO YL[0] VLO VLO VLO VLO S1AHSF400W40_CNT_CORE_F_M4
XTOPEDGE VDDHD VDD VSS WLP_SAE WLP_SAE_TK S1AHSF400W40_TOP_EDGE
XMIO_HD0 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD1 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD2 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD3 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD4 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD5 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD6 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD7 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD8 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD9 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD10 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD11 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD12 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD13 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD14 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD15 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD16 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD17 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD18 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD19 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD20 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD21 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD22 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD23 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD24 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD25 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD26 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD27 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD28 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD29 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD30 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD31 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD32 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD33 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD34 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD35 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD36 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD37 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD38 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD39 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD40 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD41 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD42 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD43 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD44 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD45 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD46 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD47 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD48 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD49 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD50 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD51 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD52 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD53 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD54 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
XMIO_HD55 VDDHD PD_BUF VDD VDD S1AHSF400W40_MIO_HD
D_WEB VSS WEB NDIO 0.056P
D_CEB VSS CEB NDIO 0.056P
D_WTESL_2 VSS WTSEL[2] NDIO 0.056P
D_WTESL_1 VSS WTSEL[1] NDIO 0.056P
D_WTESL_0 VSS WTSEL[0] NDIO 0.056P
D_RTESL_1 VSS RTSEL[1] NDIO 0.056P
D_RTESL_0 VSS RTSEL[0] NDIO 0.056P
D_CLK VSS CLK NDIO 0.056P
D_A0 VSS A[0] NDIO 0.056P
D_A1 VSS A[1] NDIO 0.056P
D_A2 VSS A[2] NDIO 0.056P
D_A3 VSS A[3] NDIO 0.056P
D_A4 VSS A[4] NDIO 0.056P
D_A5 VSS A[5] NDIO 0.056P
D_A6 VSS A[6] NDIO 0.056P
D_A7 VSS A[7] NDIO 0.056P
D_A8 VSS A[8] NDIO 0.056P
D_A9 VSS A[9] NDIO 0.056P
D_D0 VSS D[0] NDIO 0.056P
D_D1 VSS D[1] NDIO 0.056P
D_D2 VSS D[2] NDIO 0.056P
D_D3 VSS D[3] NDIO 0.056P
D_D4 VSS D[4] NDIO 0.056P
D_D5 VSS D[5] NDIO 0.056P
D_D6 VSS D[6] NDIO 0.056P
D_D7 VSS D[7] NDIO 0.056P
D_D8 VSS D[8] NDIO 0.056P
D_D9 VSS D[9] NDIO 0.056P
D_D10 VSS D[10] NDIO 0.056P
D_D11 VSS D[11] NDIO 0.056P
D_D12 VSS D[12] NDIO 0.056P
D_D13 VSS D[13] NDIO 0.056P
D_D14 VSS D[14] NDIO 0.056P
D_D15 VSS D[15] NDIO 0.056P
D_D16 VSS D[16] NDIO 0.056P
D_D17 VSS D[17] NDIO 0.056P
D_D18 VSS D[18] NDIO 0.056P
D_D19 VSS D[19] NDIO 0.056P
D_D20 VSS D[20] NDIO 0.056P
D_D21 VSS D[21] NDIO 0.056P
D_D22 VSS D[22] NDIO 0.056P
D_D23 VSS D[23] NDIO 0.056P
D_D24 VSS D[24] NDIO 0.056P
D_D25 VSS D[25] NDIO 0.056P
D_D26 VSS D[26] NDIO 0.056P
D_D27 VSS D[27] NDIO 0.056P
D_D28 VSS D[28] NDIO 0.056P
D_D29 VSS D[29] NDIO 0.056P
D_D30 VSS D[30] NDIO 0.056P
D_D31 VSS D[31] NDIO 0.056P
D_D32 VSS D[32] NDIO 0.056P
D_D33 VSS D[33] NDIO 0.056P
D_D34 VSS D[34] NDIO 0.056P
D_D35 VSS D[35] NDIO 0.056P
D_D36 VSS D[36] NDIO 0.056P
D_D37 VSS D[37] NDIO 0.056P
D_D38 VSS D[38] NDIO 0.056P
D_D39 VSS D[39] NDIO 0.056P
D_D40 VSS D[40] NDIO 0.056P
D_D41 VSS D[41] NDIO 0.056P
D_D42 VSS D[42] NDIO 0.056P
D_D43 VSS D[43] NDIO 0.056P
D_D44 VSS D[44] NDIO 0.056P
D_D45 VSS D[45] NDIO 0.056P
D_D46 VSS D[46] NDIO 0.056P
D_D47 VSS D[47] NDIO 0.056P
D_D48 VSS D[48] NDIO 0.056P
D_D49 VSS D[49] NDIO 0.056P
D_D50 VSS D[50] NDIO 0.056P
D_D51 VSS D[51] NDIO 0.056P
D_D52 VSS D[52] NDIO 0.056P
D_D53 VSS D[53] NDIO 0.056P
D_D54 VSS D[54] NDIO 0.056P
D_D55 VSS D[55] NDIO 0.056P
D_D56 VSS D[56] NDIO 0.056P
D_D57 VSS D[57] NDIO 0.056P
D_D58 VSS D[58] NDIO 0.056P
D_D59 VSS D[59] NDIO 0.056P
D_D60 VSS D[60] NDIO 0.056P
D_D61 VSS D[61] NDIO 0.056P
D_D62 VSS D[62] NDIO 0.056P
D_D63 VSS D[63] NDIO 0.056P
D_BWEB0 VSS BWEB[0] NDIO 0.056P
D_BWEB1 VSS BWEB[1] NDIO 0.056P
D_BWEB2 VSS BWEB[2] NDIO 0.056P
D_BWEB3 VSS BWEB[3] NDIO 0.056P
D_BWEB4 VSS BWEB[4] NDIO 0.056P
D_BWEB5 VSS BWEB[5] NDIO 0.056P
D_BWEB6 VSS BWEB[6] NDIO 0.056P
D_BWEB7 VSS BWEB[7] NDIO 0.056P
D_BWEB8 VSS BWEB[8] NDIO 0.056P
D_BWEB9 VSS BWEB[9] NDIO 0.056P
D_BWEB10 VSS BWEB[10] NDIO 0.056P
D_BWEB11 VSS BWEB[11] NDIO 0.056P
D_BWEB12 VSS BWEB[12] NDIO 0.056P
D_BWEB13 VSS BWEB[13] NDIO 0.056P
D_BWEB14 VSS BWEB[14] NDIO 0.056P
D_BWEB15 VSS BWEB[15] NDIO 0.056P
D_BWEB16 VSS BWEB[16] NDIO 0.056P
D_BWEB17 VSS BWEB[17] NDIO 0.056P
D_BWEB18 VSS BWEB[18] NDIO 0.056P
D_BWEB19 VSS BWEB[19] NDIO 0.056P
D_BWEB20 VSS BWEB[20] NDIO 0.056P
D_BWEB21 VSS BWEB[21] NDIO 0.056P
D_BWEB22 VSS BWEB[22] NDIO 0.056P
D_BWEB23 VSS BWEB[23] NDIO 0.056P
D_BWEB24 VSS BWEB[24] NDIO 0.056P
D_BWEB25 VSS BWEB[25] NDIO 0.056P
D_BWEB26 VSS BWEB[26] NDIO 0.056P
D_BWEB27 VSS BWEB[27] NDIO 0.056P
D_BWEB28 VSS BWEB[28] NDIO 0.056P
D_BWEB29 VSS BWEB[29] NDIO 0.056P
D_BWEB30 VSS BWEB[30] NDIO 0.056P
D_BWEB31 VSS BWEB[31] NDIO 0.056P
D_BWEB32 VSS BWEB[32] NDIO 0.056P
D_BWEB33 VSS BWEB[33] NDIO 0.056P
D_BWEB34 VSS BWEB[34] NDIO 0.056P
D_BWEB35 VSS BWEB[35] NDIO 0.056P
D_BWEB36 VSS BWEB[36] NDIO 0.056P
D_BWEB37 VSS BWEB[37] NDIO 0.056P
D_BWEB38 VSS BWEB[38] NDIO 0.056P
D_BWEB39 VSS BWEB[39] NDIO 0.056P
D_BWEB40 VSS BWEB[40] NDIO 0.056P
D_BWEB41 VSS BWEB[41] NDIO 0.056P
D_BWEB42 VSS BWEB[42] NDIO 0.056P
D_BWEB43 VSS BWEB[43] NDIO 0.056P
D_BWEB44 VSS BWEB[44] NDIO 0.056P
D_BWEB45 VSS BWEB[45] NDIO 0.056P
D_BWEB46 VSS BWEB[46] NDIO 0.056P
D_BWEB47 VSS BWEB[47] NDIO 0.056P
D_BWEB48 VSS BWEB[48] NDIO 0.056P
D_BWEB49 VSS BWEB[49] NDIO 0.056P
D_BWEB50 VSS BWEB[50] NDIO 0.056P
D_BWEB51 VSS BWEB[51] NDIO 0.056P
D_BWEB52 VSS BWEB[52] NDIO 0.056P
D_BWEB53 VSS BWEB[53] NDIO 0.056P
D_BWEB54 VSS BWEB[54] NDIO 0.056P
D_BWEB55 VSS BWEB[55] NDIO 0.056P
D_BWEB56 VSS BWEB[56] NDIO 0.056P
D_BWEB57 VSS BWEB[57] NDIO 0.056P
D_BWEB58 VSS BWEB[58] NDIO 0.056P
D_BWEB59 VSS BWEB[59] NDIO 0.056P
D_BWEB60 VSS BWEB[60] NDIO 0.056P
D_BWEB61 VSS BWEB[61] NDIO 0.056P
D_BWEB62 VSS BWEB[62] NDIO 0.056P
D_BWEB63 VSS BWEB[63] NDIO 0.056P
.ENDS

