# Created by MC2 : Version 2010.02.00.a on 2022/02/24, 21:11:02

###############################################################################
#        Software       : TSMC MEMORY COMPILER 2010.02.00.a
#        Technology     : 65 nm CMOS LOGIC Low Power LowK Cu 1P10M 1.1
#                         Standard-vt logic, cell implant SRAM bit cell
#        Memory Type    : TSMC 65nm Low Power SPHS SRAM Without Redundancy
#        Library Name   : ts1n65lphsa1024x64m4f
#        Library Version: 210a
#        Generated Time : 2022/02/24, 21:11:02
###############################################################################
#
#STATEMENT OF USE
#
#This information contains confidential and proprietary information of TSMC.
#No part of this information may be reproduced, transmitted, transcribed,
#stored in a retrieval system, or translated into any human or computer
#language, in any form or by any means, electronic, mechanical, magnetic,
#optical, chemical, manual, or otherwise, without the prior written permission
#of TSMC. This information was prepared for informational purpose and is for
#use by TSMC's customers only. TSMC reserves the right to make changes in the
#information at any time and without notice.
#
###############################################################################
 
MACRO TS1N65LPHSA1024X64M4F
	CLASS BLOCK ;
	FOREIGN TS1N65LPHSA1024X64M4F 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 306.880 BY 213.850 ;
	SYMMETRY X Y R90 ;

	PIN A[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 157.670 0.000 158.070 0.430 ;
			LAYER M1 ;
			RECT 157.670 0.000 158.070 0.430 ;
			LAYER M3 ;
			RECT 157.670 0.000 158.070 0.430 ;
		END
	END A[0]

	PIN A[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 161.430 0.000 161.830 0.430 ;
			LAYER M1 ;
			RECT 161.430 0.000 161.830 0.430 ;
			LAYER M3 ;
			RECT 161.430 0.000 161.830 0.430 ;
		END
	END A[1]

	PIN A[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 138.170 0.000 138.570 0.430 ;
			LAYER M3 ;
			RECT 138.170 0.000 138.570 0.430 ;
			LAYER M2 ;
			RECT 138.170 0.000 138.570 0.430 ;
		END
	END A[2]

	PIN A[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 141.930 0.000 142.330 0.430 ;
			LAYER M2 ;
			RECT 141.930 0.000 142.330 0.430 ;
			LAYER M3 ;
			RECT 141.930 0.000 142.330 0.430 ;
		END
	END A[3]

	PIN A[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 138.870 0.000 139.270 0.430 ;
			LAYER M2 ;
			RECT 138.870 0.000 139.270 0.430 ;
			LAYER M1 ;
			RECT 138.870 0.000 139.270 0.430 ;
		END
	END A[4]

	PIN A[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 142.630 0.000 143.030 0.430 ;
			LAYER M1 ;
			RECT 142.630 0.000 143.030 0.430 ;
			LAYER M2 ;
			RECT 142.630 0.000 143.030 0.430 ;
		END
	END A[5]

	PIN A[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 146.390 0.000 146.790 0.430 ;
			LAYER M1 ;
			RECT 146.390 0.000 146.790 0.430 ;
			LAYER M3 ;
			RECT 146.390 0.000 146.790 0.430 ;
		END
	END A[6]

	PIN A[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 145.690 0.000 146.090 0.430 ;
			LAYER M2 ;
			RECT 145.690 0.000 146.090 0.430 ;
			LAYER M3 ;
			RECT 145.690 0.000 146.090 0.430 ;
		END
	END A[7]

	PIN A[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 153.210 0.000 153.610 0.430 ;
			LAYER M3 ;
			RECT 153.210 0.000 153.610 0.430 ;
			LAYER M2 ;
			RECT 153.210 0.000 153.610 0.430 ;
		END
	END A[8]

	PIN A[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 156.970 0.000 157.370 0.430 ;
			LAYER M1 ;
			RECT 156.970 0.000 157.370 0.430 ;
			LAYER M2 ;
			RECT 156.970 0.000 157.370 0.430 ;
		END
	END A[9]

	PIN BWEB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 2.340 0.000 2.740 0.430 ;
			LAYER M1 ;
			RECT 2.340 0.000 2.740 0.430 ;
			LAYER M3 ;
			RECT 2.340 0.000 2.740 0.430 ;
		END
	END BWEB[0]

	PIN BWEB[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 44.340 0.000 44.740 0.430 ;
			LAYER M2 ;
			RECT 44.340 0.000 44.740 0.430 ;
			LAYER M3 ;
			RECT 44.340 0.000 44.740 0.430 ;
		END
	END BWEB[10]

	PIN BWEB[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 48.540 0.000 48.940 0.430 ;
			LAYER M1 ;
			RECT 48.540 0.000 48.940 0.430 ;
			LAYER M3 ;
			RECT 48.540 0.000 48.940 0.430 ;
		END
	END BWEB[11]

	PIN BWEB[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 52.740 0.000 53.140 0.430 ;
			LAYER M3 ;
			RECT 52.740 0.000 53.140 0.430 ;
			LAYER M1 ;
			RECT 52.740 0.000 53.140 0.430 ;
		END
	END BWEB[12]

	PIN BWEB[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 56.940 0.000 57.340 0.430 ;
			LAYER M3 ;
			RECT 56.940 0.000 57.340 0.430 ;
			LAYER M1 ;
			RECT 56.940 0.000 57.340 0.430 ;
		END
	END BWEB[13]

	PIN BWEB[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 61.140 0.000 61.540 0.430 ;
			LAYER M1 ;
			RECT 61.140 0.000 61.540 0.430 ;
			LAYER M3 ;
			RECT 61.140 0.000 61.540 0.430 ;
		END
	END BWEB[14]

	PIN BWEB[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 65.340 0.000 65.740 0.430 ;
			LAYER M1 ;
			RECT 65.340 0.000 65.740 0.430 ;
			LAYER M2 ;
			RECT 65.340 0.000 65.740 0.430 ;
		END
	END BWEB[15]

	PIN BWEB[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 69.540 0.000 69.940 0.430 ;
			LAYER M1 ;
			RECT 69.540 0.000 69.940 0.430 ;
			LAYER M2 ;
			RECT 69.540 0.000 69.940 0.430 ;
		END
	END BWEB[16]

	PIN BWEB[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 73.740 0.000 74.140 0.430 ;
			LAYER M3 ;
			RECT 73.740 0.000 74.140 0.430 ;
			LAYER M1 ;
			RECT 73.740 0.000 74.140 0.430 ;
		END
	END BWEB[17]

	PIN BWEB[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 77.940 0.000 78.340 0.430 ;
			LAYER M3 ;
			RECT 77.940 0.000 78.340 0.430 ;
			LAYER M1 ;
			RECT 77.940 0.000 78.340 0.430 ;
		END
	END BWEB[18]

	PIN BWEB[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 82.140 0.000 82.540 0.430 ;
			LAYER M2 ;
			RECT 82.140 0.000 82.540 0.430 ;
			LAYER M3 ;
			RECT 82.140 0.000 82.540 0.430 ;
		END
	END BWEB[19]

	PIN BWEB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 6.540 0.000 6.940 0.430 ;
			LAYER M1 ;
			RECT 6.540 0.000 6.940 0.430 ;
			LAYER M3 ;
			RECT 6.540 0.000 6.940 0.430 ;
		END
	END BWEB[1]

	PIN BWEB[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 86.340 0.000 86.740 0.430 ;
			LAYER M1 ;
			RECT 86.340 0.000 86.740 0.430 ;
			LAYER M2 ;
			RECT 86.340 0.000 86.740 0.430 ;
		END
	END BWEB[20]

	PIN BWEB[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 90.540 0.000 90.940 0.430 ;
			LAYER M3 ;
			RECT 90.540 0.000 90.940 0.430 ;
			LAYER M1 ;
			RECT 90.540 0.000 90.940 0.430 ;
		END
	END BWEB[21]

	PIN BWEB[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 94.740 0.000 95.140 0.430 ;
			LAYER M1 ;
			RECT 94.740 0.000 95.140 0.430 ;
			LAYER M2 ;
			RECT 94.740 0.000 95.140 0.430 ;
		END
	END BWEB[22]

	PIN BWEB[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 98.940 0.000 99.340 0.430 ;
			LAYER M1 ;
			RECT 98.940 0.000 99.340 0.430 ;
			LAYER M2 ;
			RECT 98.940 0.000 99.340 0.430 ;
		END
	END BWEB[23]

	PIN BWEB[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 103.140 0.000 103.540 0.430 ;
			LAYER M1 ;
			RECT 103.140 0.000 103.540 0.430 ;
			LAYER M3 ;
			RECT 103.140 0.000 103.540 0.430 ;
		END
	END BWEB[24]

	PIN BWEB[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 107.340 0.000 107.740 0.430 ;
			LAYER M1 ;
			RECT 107.340 0.000 107.740 0.430 ;
			LAYER M3 ;
			RECT 107.340 0.000 107.740 0.430 ;
		END
	END BWEB[25]

	PIN BWEB[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 111.540 0.000 111.940 0.430 ;
			LAYER M1 ;
			RECT 111.540 0.000 111.940 0.430 ;
			LAYER M2 ;
			RECT 111.540 0.000 111.940 0.430 ;
		END
	END BWEB[26]

	PIN BWEB[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 115.740 0.000 116.140 0.430 ;
			LAYER M1 ;
			RECT 115.740 0.000 116.140 0.430 ;
			LAYER M3 ;
			RECT 115.740 0.000 116.140 0.430 ;
		END
	END BWEB[27]

	PIN BWEB[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 119.630 0.000 120.030 0.430 ;
			LAYER M1 ;
			RECT 119.630 0.000 120.030 0.430 ;
			LAYER M2 ;
			RECT 119.630 0.000 120.030 0.430 ;
		END
	END BWEB[28]

	PIN BWEB[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 123.820 0.000 124.220 0.430 ;
			LAYER M3 ;
			RECT 123.820 0.000 124.220 0.430 ;
			LAYER M2 ;
			RECT 123.820 0.000 124.220 0.430 ;
		END
	END BWEB[29]

	PIN BWEB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 10.740 0.000 11.140 0.430 ;
			LAYER M2 ;
			RECT 10.740 0.000 11.140 0.430 ;
			LAYER M1 ;
			RECT 10.740 0.000 11.140 0.430 ;
		END
	END BWEB[2]

	PIN BWEB[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 127.650 0.000 128.050 0.430 ;
			LAYER M3 ;
			RECT 127.650 0.000 128.050 0.430 ;
			LAYER M1 ;
			RECT 127.650 0.000 128.050 0.430 ;
		END
	END BWEB[30]

	PIN BWEB[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 131.880 0.000 132.280 0.430 ;
			LAYER M2 ;
			RECT 131.880 0.000 132.280 0.430 ;
			LAYER M3 ;
			RECT 131.880 0.000 132.280 0.430 ;
		END
	END BWEB[31]

	PIN BWEB[32]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 171.645 0.000 172.045 0.430 ;
			LAYER M2 ;
			RECT 171.645 0.000 172.045 0.430 ;
			LAYER M3 ;
			RECT 171.645 0.000 172.045 0.430 ;
		END
	END BWEB[32]

	PIN BWEB[33]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 175.895 0.000 176.295 0.430 ;
			LAYER M1 ;
			RECT 175.895 0.000 176.295 0.430 ;
			LAYER M3 ;
			RECT 175.895 0.000 176.295 0.430 ;
		END
	END BWEB[33]

	PIN BWEB[34]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 179.905 0.000 180.305 0.430 ;
			LAYER M1 ;
			RECT 179.905 0.000 180.305 0.430 ;
			LAYER M2 ;
			RECT 179.905 0.000 180.305 0.430 ;
		END
	END BWEB[34]

	PIN BWEB[35]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 183.395 0.000 183.795 0.430 ;
			LAYER M3 ;
			RECT 183.395 0.000 183.795 0.430 ;
			LAYER M2 ;
			RECT 183.395 0.000 183.795 0.430 ;
		END
	END BWEB[35]

	PIN BWEB[36]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 188.340 0.000 188.740 0.430 ;
			LAYER M3 ;
			RECT 188.340 0.000 188.740 0.430 ;
			LAYER M1 ;
			RECT 188.340 0.000 188.740 0.430 ;
		END
	END BWEB[36]

	PIN BWEB[37]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 192.540 0.000 192.940 0.430 ;
			LAYER M2 ;
			RECT 192.540 0.000 192.940 0.430 ;
			LAYER M3 ;
			RECT 192.540 0.000 192.940 0.430 ;
		END
	END BWEB[37]

	PIN BWEB[38]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 196.740 0.000 197.140 0.430 ;
			LAYER M3 ;
			RECT 196.740 0.000 197.140 0.430 ;
			LAYER M2 ;
			RECT 196.740 0.000 197.140 0.430 ;
		END
	END BWEB[38]

	PIN BWEB[39]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 200.940 0.000 201.340 0.430 ;
			LAYER M3 ;
			RECT 200.940 0.000 201.340 0.430 ;
			LAYER M1 ;
			RECT 200.940 0.000 201.340 0.430 ;
		END
	END BWEB[39]

	PIN BWEB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 14.940 0.000 15.340 0.430 ;
			LAYER M3 ;
			RECT 14.940 0.000 15.340 0.430 ;
			LAYER M1 ;
			RECT 14.940 0.000 15.340 0.430 ;
		END
	END BWEB[3]

	PIN BWEB[40]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 205.140 0.000 205.540 0.430 ;
			LAYER M2 ;
			RECT 205.140 0.000 205.540 0.430 ;
			LAYER M3 ;
			RECT 205.140 0.000 205.540 0.430 ;
		END
	END BWEB[40]

	PIN BWEB[41]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 209.340 0.000 209.740 0.430 ;
			LAYER M1 ;
			RECT 209.340 0.000 209.740 0.430 ;
			LAYER M2 ;
			RECT 209.340 0.000 209.740 0.430 ;
		END
	END BWEB[41]

	PIN BWEB[42]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 213.540 0.000 213.940 0.430 ;
			LAYER M3 ;
			RECT 213.540 0.000 213.940 0.430 ;
			LAYER M1 ;
			RECT 213.540 0.000 213.940 0.430 ;
		END
	END BWEB[42]

	PIN BWEB[43]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 217.740 0.000 218.140 0.430 ;
			LAYER M1 ;
			RECT 217.740 0.000 218.140 0.430 ;
			LAYER M2 ;
			RECT 217.740 0.000 218.140 0.430 ;
		END
	END BWEB[43]

	PIN BWEB[44]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 221.940 0.000 222.340 0.430 ;
			LAYER M3 ;
			RECT 221.940 0.000 222.340 0.430 ;
			LAYER M1 ;
			RECT 221.940 0.000 222.340 0.430 ;
		END
	END BWEB[44]

	PIN BWEB[45]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 226.140 0.000 226.540 0.430 ;
			LAYER M3 ;
			RECT 226.140 0.000 226.540 0.430 ;
			LAYER M2 ;
			RECT 226.140 0.000 226.540 0.430 ;
		END
	END BWEB[45]

	PIN BWEB[46]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 230.340 0.000 230.740 0.430 ;
			LAYER M1 ;
			RECT 230.340 0.000 230.740 0.430 ;
			LAYER M2 ;
			RECT 230.340 0.000 230.740 0.430 ;
		END
	END BWEB[46]

	PIN BWEB[47]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 234.540 0.000 234.940 0.430 ;
			LAYER M3 ;
			RECT 234.540 0.000 234.940 0.430 ;
			LAYER M2 ;
			RECT 234.540 0.000 234.940 0.430 ;
		END
	END BWEB[47]

	PIN BWEB[48]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 238.740 0.000 239.140 0.430 ;
			LAYER M3 ;
			RECT 238.740 0.000 239.140 0.430 ;
			LAYER M1 ;
			RECT 238.740 0.000 239.140 0.430 ;
		END
	END BWEB[48]

	PIN BWEB[49]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 242.940 0.000 243.340 0.430 ;
			LAYER M3 ;
			RECT 242.940 0.000 243.340 0.430 ;
			LAYER M2 ;
			RECT 242.940 0.000 243.340 0.430 ;
		END
	END BWEB[49]

	PIN BWEB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 19.140 0.000 19.540 0.430 ;
			LAYER M1 ;
			RECT 19.140 0.000 19.540 0.430 ;
			LAYER M2 ;
			RECT 19.140 0.000 19.540 0.430 ;
		END
	END BWEB[4]

	PIN BWEB[50]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 247.140 0.000 247.540 0.430 ;
			LAYER M3 ;
			RECT 247.140 0.000 247.540 0.430 ;
			LAYER M1 ;
			RECT 247.140 0.000 247.540 0.430 ;
		END
	END BWEB[50]

	PIN BWEB[51]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 251.340 0.000 251.740 0.430 ;
			LAYER M2 ;
			RECT 251.340 0.000 251.740 0.430 ;
			LAYER M3 ;
			RECT 251.340 0.000 251.740 0.430 ;
		END
	END BWEB[51]

	PIN BWEB[52]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 255.540 0.000 255.940 0.430 ;
			LAYER M2 ;
			RECT 255.540 0.000 255.940 0.430 ;
			LAYER M3 ;
			RECT 255.540 0.000 255.940 0.430 ;
		END
	END BWEB[52]

	PIN BWEB[53]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 259.740 0.000 260.140 0.430 ;
			LAYER M3 ;
			RECT 259.740 0.000 260.140 0.430 ;
			LAYER M1 ;
			RECT 259.740 0.000 260.140 0.430 ;
		END
	END BWEB[53]

	PIN BWEB[54]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 263.940 0.000 264.340 0.430 ;
			LAYER M1 ;
			RECT 263.940 0.000 264.340 0.430 ;
			LAYER M2 ;
			RECT 263.940 0.000 264.340 0.430 ;
		END
	END BWEB[54]

	PIN BWEB[55]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 268.140 0.000 268.540 0.430 ;
			LAYER M3 ;
			RECT 268.140 0.000 268.540 0.430 ;
			LAYER M2 ;
			RECT 268.140 0.000 268.540 0.430 ;
		END
	END BWEB[55]

	PIN BWEB[56]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 272.340 0.000 272.740 0.430 ;
			LAYER M1 ;
			RECT 272.340 0.000 272.740 0.430 ;
			LAYER M3 ;
			RECT 272.340 0.000 272.740 0.430 ;
		END
	END BWEB[56]

	PIN BWEB[57]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 276.540 0.000 276.940 0.430 ;
			LAYER M3 ;
			RECT 276.540 0.000 276.940 0.430 ;
			LAYER M1 ;
			RECT 276.540 0.000 276.940 0.430 ;
		END
	END BWEB[57]

	PIN BWEB[58]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 280.740 0.000 281.140 0.430 ;
			LAYER M3 ;
			RECT 280.740 0.000 281.140 0.430 ;
			LAYER M1 ;
			RECT 280.740 0.000 281.140 0.430 ;
		END
	END BWEB[58]

	PIN BWEB[59]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 284.940 0.000 285.340 0.430 ;
			LAYER M3 ;
			RECT 284.940 0.000 285.340 0.430 ;
			LAYER M1 ;
			RECT 284.940 0.000 285.340 0.430 ;
		END
	END BWEB[59]

	PIN BWEB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 23.340 0.000 23.740 0.430 ;
			LAYER M2 ;
			RECT 23.340 0.000 23.740 0.430 ;
			LAYER M1 ;
			RECT 23.340 0.000 23.740 0.430 ;
		END
	END BWEB[5]

	PIN BWEB[60]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 289.140 0.000 289.540 0.430 ;
			LAYER M1 ;
			RECT 289.140 0.000 289.540 0.430 ;
			LAYER M2 ;
			RECT 289.140 0.000 289.540 0.430 ;
		END
	END BWEB[60]

	PIN BWEB[61]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 293.340 0.000 293.740 0.430 ;
			LAYER M2 ;
			RECT 293.340 0.000 293.740 0.430 ;
			LAYER M3 ;
			RECT 293.340 0.000 293.740 0.430 ;
		END
	END BWEB[61]

	PIN BWEB[62]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 297.540 0.000 297.940 0.430 ;
			LAYER M2 ;
			RECT 297.540 0.000 297.940 0.430 ;
			LAYER M3 ;
			RECT 297.540 0.000 297.940 0.430 ;
		END
	END BWEB[62]

	PIN BWEB[63]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 301.740 0.000 302.140 0.430 ;
			LAYER M2 ;
			RECT 301.740 0.000 302.140 0.430 ;
			LAYER M3 ;
			RECT 301.740 0.000 302.140 0.430 ;
		END
	END BWEB[63]

	PIN BWEB[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 27.540 0.000 27.940 0.430 ;
			LAYER M1 ;
			RECT 27.540 0.000 27.940 0.430 ;
			LAYER M2 ;
			RECT 27.540 0.000 27.940 0.430 ;
		END
	END BWEB[6]

	PIN BWEB[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 31.740 0.000 32.140 0.430 ;
			LAYER M1 ;
			RECT 31.740 0.000 32.140 0.430 ;
			LAYER M3 ;
			RECT 31.740 0.000 32.140 0.430 ;
		END
	END BWEB[7]

	PIN BWEB[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 35.940 0.000 36.340 0.430 ;
			LAYER M2 ;
			RECT 35.940 0.000 36.340 0.430 ;
			LAYER M3 ;
			RECT 35.940 0.000 36.340 0.430 ;
		END
	END BWEB[8]

	PIN BWEB[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 40.140 0.000 40.540 0.430 ;
			LAYER M1 ;
			RECT 40.140 0.000 40.540 0.430 ;
			LAYER M2 ;
			RECT 40.140 0.000 40.540 0.430 ;
		END
	END BWEB[9]

	PIN CEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 169.580 0.000 169.980 0.430 ;
			LAYER M1 ;
			RECT 169.580 0.000 169.980 0.430 ;
			LAYER M2 ;
			RECT 169.580 0.000 169.980 0.430 ;
		END
	END CEB

	PIN CLK
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 167.270 0.000 167.670 0.430 ;
			LAYER M3 ;
			RECT 167.270 0.000 167.670 0.430 ;
			LAYER M2 ;
			RECT 167.270 0.000 167.670 0.430 ;
		END
	END CLK

	PIN D[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 4.740 0.000 5.140 0.430 ;
			LAYER M3 ;
			RECT 4.740 0.000 5.140 0.430 ;
			LAYER M1 ;
			RECT 4.740 0.000 5.140 0.430 ;
		END
	END D[0]

	PIN D[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 46.740 0.000 47.140 0.430 ;
			LAYER M2 ;
			RECT 46.740 0.000 47.140 0.430 ;
			LAYER M1 ;
			RECT 46.740 0.000 47.140 0.430 ;
		END
	END D[10]

	PIN D[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 50.940 0.000 51.340 0.430 ;
			LAYER M2 ;
			RECT 50.940 0.000 51.340 0.430 ;
			LAYER M3 ;
			RECT 50.940 0.000 51.340 0.430 ;
		END
	END D[11]

	PIN D[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 55.140 0.000 55.540 0.430 ;
			LAYER M2 ;
			RECT 55.140 0.000 55.540 0.430 ;
			LAYER M3 ;
			RECT 55.140 0.000 55.540 0.430 ;
		END
	END D[12]

	PIN D[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 59.340 0.000 59.740 0.430 ;
			LAYER M3 ;
			RECT 59.340 0.000 59.740 0.430 ;
			LAYER M1 ;
			RECT 59.340 0.000 59.740 0.430 ;
		END
	END D[13]

	PIN D[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 63.540 0.000 63.940 0.430 ;
			LAYER M2 ;
			RECT 63.540 0.000 63.940 0.430 ;
			LAYER M3 ;
			RECT 63.540 0.000 63.940 0.430 ;
		END
	END D[14]

	PIN D[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 67.740 0.000 68.140 0.430 ;
			LAYER M2 ;
			RECT 67.740 0.000 68.140 0.430 ;
			LAYER M3 ;
			RECT 67.740 0.000 68.140 0.430 ;
		END
	END D[15]

	PIN D[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 71.940 0.000 72.340 0.430 ;
			LAYER M1 ;
			RECT 71.940 0.000 72.340 0.430 ;
			LAYER M2 ;
			RECT 71.940 0.000 72.340 0.430 ;
		END
	END D[16]

	PIN D[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 76.140 0.000 76.540 0.430 ;
			LAYER M1 ;
			RECT 76.140 0.000 76.540 0.430 ;
			LAYER M2 ;
			RECT 76.140 0.000 76.540 0.430 ;
		END
	END D[17]

	PIN D[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 80.340 0.000 80.740 0.430 ;
			LAYER M3 ;
			RECT 80.340 0.000 80.740 0.430 ;
			LAYER M1 ;
			RECT 80.340 0.000 80.740 0.430 ;
		END
	END D[18]

	PIN D[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 84.540 0.000 84.940 0.430 ;
			LAYER M3 ;
			RECT 84.540 0.000 84.940 0.430 ;
			LAYER M1 ;
			RECT 84.540 0.000 84.940 0.430 ;
		END
	END D[19]

	PIN D[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 8.940 0.000 9.340 0.430 ;
			LAYER M3 ;
			RECT 8.940 0.000 9.340 0.430 ;
			LAYER M1 ;
			RECT 8.940 0.000 9.340 0.430 ;
		END
	END D[1]

	PIN D[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 88.740 0.000 89.140 0.430 ;
			LAYER M3 ;
			RECT 88.740 0.000 89.140 0.430 ;
			LAYER M1 ;
			RECT 88.740 0.000 89.140 0.430 ;
		END
	END D[20]

	PIN D[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 92.940 0.000 93.340 0.430 ;
			LAYER M3 ;
			RECT 92.940 0.000 93.340 0.430 ;
			LAYER M1 ;
			RECT 92.940 0.000 93.340 0.430 ;
		END
	END D[21]

	PIN D[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 97.140 0.000 97.540 0.430 ;
			LAYER M1 ;
			RECT 97.140 0.000 97.540 0.430 ;
			LAYER M3 ;
			RECT 97.140 0.000 97.540 0.430 ;
		END
	END D[22]

	PIN D[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 101.340 0.000 101.740 0.430 ;
			LAYER M1 ;
			RECT 101.340 0.000 101.740 0.430 ;
			LAYER M3 ;
			RECT 101.340 0.000 101.740 0.430 ;
		END
	END D[23]

	PIN D[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 105.540 0.000 105.940 0.430 ;
			LAYER M1 ;
			RECT 105.540 0.000 105.940 0.430 ;
			LAYER M2 ;
			RECT 105.540 0.000 105.940 0.430 ;
		END
	END D[24]

	PIN D[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 109.740 0.000 110.140 0.430 ;
			LAYER M2 ;
			RECT 109.740 0.000 110.140 0.430 ;
			LAYER M3 ;
			RECT 109.740 0.000 110.140 0.430 ;
		END
	END D[25]

	PIN D[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 113.940 0.000 114.340 0.430 ;
			LAYER M2 ;
			RECT 113.940 0.000 114.340 0.430 ;
			LAYER M3 ;
			RECT 113.940 0.000 114.340 0.430 ;
		END
	END D[26]

	PIN D[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 118.140 0.000 118.540 0.430 ;
			LAYER M2 ;
			RECT 118.140 0.000 118.540 0.430 ;
			LAYER M3 ;
			RECT 118.140 0.000 118.540 0.430 ;
		END
	END D[27]

	PIN D[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 122.710 0.000 123.110 0.430 ;
			LAYER M3 ;
			RECT 122.710 0.000 123.110 0.430 ;
			LAYER M1 ;
			RECT 122.710 0.000 123.110 0.430 ;
		END
	END D[28]

	PIN D[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 126.980 0.000 127.380 0.430 ;
			LAYER M3 ;
			RECT 126.980 0.000 127.380 0.430 ;
			LAYER M1 ;
			RECT 126.980 0.000 127.380 0.430 ;
		END
	END D[29]

	PIN D[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 13.140 0.000 13.540 0.430 ;
			LAYER M1 ;
			RECT 13.140 0.000 13.540 0.430 ;
			LAYER M3 ;
			RECT 13.140 0.000 13.540 0.430 ;
		END
	END D[2]

	PIN D[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 130.670 0.000 131.070 0.430 ;
			LAYER M1 ;
			RECT 130.670 0.000 131.070 0.430 ;
			LAYER M3 ;
			RECT 130.670 0.000 131.070 0.430 ;
		END
	END D[30]

	PIN D[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 135.160 0.000 135.560 0.430 ;
			LAYER M1 ;
			RECT 135.160 0.000 135.560 0.430 ;
			LAYER M3 ;
			RECT 135.160 0.000 135.560 0.430 ;
		END
	END D[31]

	PIN D[32]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 174.645 0.000 175.045 0.430 ;
			LAYER M3 ;
			RECT 174.645 0.000 175.045 0.430 ;
			LAYER M1 ;
			RECT 174.645 0.000 175.045 0.430 ;
		END
	END D[32]

	PIN D[33]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 178.615 0.000 179.015 0.430 ;
			LAYER M3 ;
			RECT 178.615 0.000 179.015 0.430 ;
			LAYER M1 ;
			RECT 178.615 0.000 179.015 0.430 ;
		END
	END D[33]

	PIN D[34]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 182.795 0.000 183.195 0.430 ;
			LAYER M3 ;
			RECT 182.795 0.000 183.195 0.430 ;
			LAYER M2 ;
			RECT 182.795 0.000 183.195 0.430 ;
		END
	END D[34]

	PIN D[35]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 187.050 0.000 187.450 0.430 ;
			LAYER M2 ;
			RECT 187.050 0.000 187.450 0.430 ;
			LAYER M1 ;
			RECT 187.050 0.000 187.450 0.430 ;
		END
	END D[35]

	PIN D[36]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 190.740 0.000 191.140 0.430 ;
			LAYER M3 ;
			RECT 190.740 0.000 191.140 0.430 ;
			LAYER M1 ;
			RECT 190.740 0.000 191.140 0.430 ;
		END
	END D[36]

	PIN D[37]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 194.940 0.000 195.340 0.430 ;
			LAYER M3 ;
			RECT 194.940 0.000 195.340 0.430 ;
			LAYER M1 ;
			RECT 194.940 0.000 195.340 0.430 ;
		END
	END D[37]

	PIN D[38]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 199.140 0.000 199.540 0.430 ;
			LAYER M3 ;
			RECT 199.140 0.000 199.540 0.430 ;
			LAYER M1 ;
			RECT 199.140 0.000 199.540 0.430 ;
		END
	END D[38]

	PIN D[39]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 203.340 0.000 203.740 0.430 ;
			LAYER M1 ;
			RECT 203.340 0.000 203.740 0.430 ;
			LAYER M2 ;
			RECT 203.340 0.000 203.740 0.430 ;
		END
	END D[39]

	PIN D[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.340 0.000 17.740 0.430 ;
			LAYER M2 ;
			RECT 17.340 0.000 17.740 0.430 ;
			LAYER M3 ;
			RECT 17.340 0.000 17.740 0.430 ;
		END
	END D[3]

	PIN D[40]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 207.540 0.000 207.940 0.430 ;
			LAYER M2 ;
			RECT 207.540 0.000 207.940 0.430 ;
			LAYER M1 ;
			RECT 207.540 0.000 207.940 0.430 ;
		END
	END D[40]

	PIN D[41]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 211.740 0.000 212.140 0.430 ;
			LAYER M3 ;
			RECT 211.740 0.000 212.140 0.430 ;
			LAYER M1 ;
			RECT 211.740 0.000 212.140 0.430 ;
		END
	END D[41]

	PIN D[42]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 215.940 0.000 216.340 0.430 ;
			LAYER M2 ;
			RECT 215.940 0.000 216.340 0.430 ;
			LAYER M3 ;
			RECT 215.940 0.000 216.340 0.430 ;
		END
	END D[42]

	PIN D[43]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 220.140 0.000 220.540 0.430 ;
			LAYER M1 ;
			RECT 220.140 0.000 220.540 0.430 ;
			LAYER M2 ;
			RECT 220.140 0.000 220.540 0.430 ;
		END
	END D[43]

	PIN D[44]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 224.340 0.000 224.740 0.430 ;
			LAYER M1 ;
			RECT 224.340 0.000 224.740 0.430 ;
			LAYER M3 ;
			RECT 224.340 0.000 224.740 0.430 ;
		END
	END D[44]

	PIN D[45]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 228.540 0.000 228.940 0.430 ;
			LAYER M1 ;
			RECT 228.540 0.000 228.940 0.430 ;
			LAYER M3 ;
			RECT 228.540 0.000 228.940 0.430 ;
		END
	END D[45]

	PIN D[46]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 232.740 0.000 233.140 0.430 ;
			LAYER M1 ;
			RECT 232.740 0.000 233.140 0.430 ;
			LAYER M3 ;
			RECT 232.740 0.000 233.140 0.430 ;
		END
	END D[46]

	PIN D[47]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 236.940 0.000 237.340 0.430 ;
			LAYER M1 ;
			RECT 236.940 0.000 237.340 0.430 ;
			LAYER M2 ;
			RECT 236.940 0.000 237.340 0.430 ;
		END
	END D[47]

	PIN D[48]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 241.140 0.000 241.540 0.430 ;
			LAYER M2 ;
			RECT 241.140 0.000 241.540 0.430 ;
			LAYER M3 ;
			RECT 241.140 0.000 241.540 0.430 ;
		END
	END D[48]

	PIN D[49]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 245.340 0.000 245.740 0.430 ;
			LAYER M2 ;
			RECT 245.340 0.000 245.740 0.430 ;
			LAYER M3 ;
			RECT 245.340 0.000 245.740 0.430 ;
		END
	END D[49]

	PIN D[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 21.540 0.000 21.940 0.430 ;
			LAYER M3 ;
			RECT 21.540 0.000 21.940 0.430 ;
			LAYER M1 ;
			RECT 21.540 0.000 21.940 0.430 ;
		END
	END D[4]

	PIN D[50]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 249.540 0.000 249.940 0.430 ;
			LAYER M1 ;
			RECT 249.540 0.000 249.940 0.430 ;
			LAYER M3 ;
			RECT 249.540 0.000 249.940 0.430 ;
		END
	END D[50]

	PIN D[51]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 253.740 0.000 254.140 0.430 ;
			LAYER M1 ;
			RECT 253.740 0.000 254.140 0.430 ;
			LAYER M2 ;
			RECT 253.740 0.000 254.140 0.430 ;
		END
	END D[51]

	PIN D[52]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 257.940 0.000 258.340 0.430 ;
			LAYER M3 ;
			RECT 257.940 0.000 258.340 0.430 ;
			LAYER M1 ;
			RECT 257.940 0.000 258.340 0.430 ;
		END
	END D[52]

	PIN D[53]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 262.140 0.000 262.540 0.430 ;
			LAYER M1 ;
			RECT 262.140 0.000 262.540 0.430 ;
			LAYER M3 ;
			RECT 262.140 0.000 262.540 0.430 ;
		END
	END D[53]

	PIN D[54]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 266.340 0.000 266.740 0.430 ;
			LAYER M3 ;
			RECT 266.340 0.000 266.740 0.430 ;
			LAYER M1 ;
			RECT 266.340 0.000 266.740 0.430 ;
		END
	END D[54]

	PIN D[55]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 270.540 0.000 270.940 0.430 ;
			LAYER M2 ;
			RECT 270.540 0.000 270.940 0.430 ;
			LAYER M3 ;
			RECT 270.540 0.000 270.940 0.430 ;
		END
	END D[55]

	PIN D[56]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 274.740 0.000 275.140 0.430 ;
			LAYER M1 ;
			RECT 274.740 0.000 275.140 0.430 ;
			LAYER M2 ;
			RECT 274.740 0.000 275.140 0.430 ;
		END
	END D[56]

	PIN D[57]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 278.940 0.000 279.340 0.430 ;
			LAYER M2 ;
			RECT 278.940 0.000 279.340 0.430 ;
			LAYER M3 ;
			RECT 278.940 0.000 279.340 0.430 ;
		END
	END D[57]

	PIN D[58]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 283.140 0.000 283.540 0.430 ;
			LAYER M3 ;
			RECT 283.140 0.000 283.540 0.430 ;
			LAYER M1 ;
			RECT 283.140 0.000 283.540 0.430 ;
		END
	END D[58]

	PIN D[59]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 287.340 0.000 287.740 0.430 ;
			LAYER M2 ;
			RECT 287.340 0.000 287.740 0.430 ;
			LAYER M3 ;
			RECT 287.340 0.000 287.740 0.430 ;
		END
	END D[59]

	PIN D[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 25.740 0.000 26.140 0.430 ;
			LAYER M1 ;
			RECT 25.740 0.000 26.140 0.430 ;
			LAYER M2 ;
			RECT 25.740 0.000 26.140 0.430 ;
		END
	END D[5]

	PIN D[60]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 291.540 0.000 291.940 0.430 ;
			LAYER M1 ;
			RECT 291.540 0.000 291.940 0.430 ;
			LAYER M2 ;
			RECT 291.540 0.000 291.940 0.430 ;
		END
	END D[60]

	PIN D[61]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 295.740 0.000 296.140 0.430 ;
			LAYER M3 ;
			RECT 295.740 0.000 296.140 0.430 ;
			LAYER M1 ;
			RECT 295.740 0.000 296.140 0.430 ;
		END
	END D[61]

	PIN D[62]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 299.940 0.000 300.340 0.430 ;
			LAYER M3 ;
			RECT 299.940 0.000 300.340 0.430 ;
			LAYER M1 ;
			RECT 299.940 0.000 300.340 0.430 ;
		END
	END D[62]

	PIN D[63]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 304.140 0.000 304.540 0.430 ;
			LAYER M2 ;
			RECT 304.140 0.000 304.540 0.430 ;
			LAYER M3 ;
			RECT 304.140 0.000 304.540 0.430 ;
		END
	END D[63]

	PIN D[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 29.940 0.000 30.340 0.430 ;
			LAYER M3 ;
			RECT 29.940 0.000 30.340 0.430 ;
			LAYER M1 ;
			RECT 29.940 0.000 30.340 0.430 ;
		END
	END D[6]

	PIN D[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 34.140 0.000 34.540 0.430 ;
			LAYER M2 ;
			RECT 34.140 0.000 34.540 0.430 ;
			LAYER M3 ;
			RECT 34.140 0.000 34.540 0.430 ;
		END
	END D[7]

	PIN D[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 38.340 0.000 38.740 0.430 ;
			LAYER M1 ;
			RECT 38.340 0.000 38.740 0.430 ;
			LAYER M2 ;
			RECT 38.340 0.000 38.740 0.430 ;
		END
	END D[8]

	PIN D[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 42.540 0.000 42.940 0.430 ;
			LAYER M1 ;
			RECT 42.540 0.000 42.940 0.430 ;
			LAYER M2 ;
			RECT 42.540 0.000 42.940 0.430 ;
		END
	END D[9]

	PIN Q[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 3.540 0.000 3.940 0.430 ;
			LAYER M3 ;
			RECT 3.540 0.000 3.940 0.430 ;
			LAYER M1 ;
			RECT 3.540 0.000 3.940 0.430 ;
		END
	END Q[0]

	PIN Q[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 45.540 0.000 45.940 0.430 ;
			LAYER M3 ;
			RECT 45.540 0.000 45.940 0.430 ;
			LAYER M2 ;
			RECT 45.540 0.000 45.940 0.430 ;
		END
	END Q[10]

	PIN Q[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 49.740 0.000 50.140 0.430 ;
			LAYER M2 ;
			RECT 49.740 0.000 50.140 0.430 ;
			LAYER M1 ;
			RECT 49.740 0.000 50.140 0.430 ;
		END
	END Q[11]

	PIN Q[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 53.940 0.000 54.340 0.430 ;
			LAYER M1 ;
			RECT 53.940 0.000 54.340 0.430 ;
			LAYER M2 ;
			RECT 53.940 0.000 54.340 0.430 ;
		END
	END Q[12]

	PIN Q[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 58.140 0.000 58.540 0.430 ;
			LAYER M2 ;
			RECT 58.140 0.000 58.540 0.430 ;
			LAYER M3 ;
			RECT 58.140 0.000 58.540 0.430 ;
		END
	END Q[13]

	PIN Q[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 62.340 0.000 62.740 0.430 ;
			LAYER M3 ;
			RECT 62.340 0.000 62.740 0.430 ;
			LAYER M2 ;
			RECT 62.340 0.000 62.740 0.430 ;
		END
	END Q[14]

	PIN Q[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 66.540 0.000 66.940 0.430 ;
			LAYER M2 ;
			RECT 66.540 0.000 66.940 0.430 ;
			LAYER M3 ;
			RECT 66.540 0.000 66.940 0.430 ;
		END
	END Q[15]

	PIN Q[16]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 70.740 0.000 71.140 0.430 ;
			LAYER M2 ;
			RECT 70.740 0.000 71.140 0.430 ;
			LAYER M1 ;
			RECT 70.740 0.000 71.140 0.430 ;
		END
	END Q[16]

	PIN Q[17]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 74.940 0.000 75.340 0.430 ;
			LAYER M3 ;
			RECT 74.940 0.000 75.340 0.430 ;
			LAYER M1 ;
			RECT 74.940 0.000 75.340 0.430 ;
		END
	END Q[17]

	PIN Q[18]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 79.140 0.000 79.540 0.430 ;
			LAYER M3 ;
			RECT 79.140 0.000 79.540 0.430 ;
			LAYER M2 ;
			RECT 79.140 0.000 79.540 0.430 ;
		END
	END Q[18]

	PIN Q[19]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 83.340 0.000 83.740 0.430 ;
			LAYER M2 ;
			RECT 83.340 0.000 83.740 0.430 ;
			LAYER M3 ;
			RECT 83.340 0.000 83.740 0.430 ;
		END
	END Q[19]

	PIN Q[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 7.740 0.000 8.140 0.430 ;
			LAYER M1 ;
			RECT 7.740 0.000 8.140 0.430 ;
			LAYER M3 ;
			RECT 7.740 0.000 8.140 0.430 ;
		END
	END Q[1]

	PIN Q[20]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 87.540 0.000 87.940 0.430 ;
			LAYER M3 ;
			RECT 87.540 0.000 87.940 0.430 ;
			LAYER M2 ;
			RECT 87.540 0.000 87.940 0.430 ;
		END
	END Q[20]

	PIN Q[21]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 91.740 0.000 92.140 0.430 ;
			LAYER M3 ;
			RECT 91.740 0.000 92.140 0.430 ;
			LAYER M2 ;
			RECT 91.740 0.000 92.140 0.430 ;
		END
	END Q[21]

	PIN Q[22]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 95.940 0.000 96.340 0.430 ;
			LAYER M2 ;
			RECT 95.940 0.000 96.340 0.430 ;
			LAYER M3 ;
			RECT 95.940 0.000 96.340 0.430 ;
		END
	END Q[22]

	PIN Q[23]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 100.140 0.000 100.540 0.430 ;
			LAYER M2 ;
			RECT 100.140 0.000 100.540 0.430 ;
			LAYER M3 ;
			RECT 100.140 0.000 100.540 0.430 ;
		END
	END Q[23]

	PIN Q[24]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 104.340 0.000 104.740 0.430 ;
			LAYER M3 ;
			RECT 104.340 0.000 104.740 0.430 ;
			LAYER M2 ;
			RECT 104.340 0.000 104.740 0.430 ;
		END
	END Q[24]

	PIN Q[25]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 108.540 0.000 108.940 0.430 ;
			LAYER M3 ;
			RECT 108.540 0.000 108.940 0.430 ;
			LAYER M2 ;
			RECT 108.540 0.000 108.940 0.430 ;
		END
	END Q[25]

	PIN Q[26]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 112.740 0.000 113.140 0.430 ;
			LAYER M3 ;
			RECT 112.740 0.000 113.140 0.430 ;
			LAYER M2 ;
			RECT 112.740 0.000 113.140 0.430 ;
		END
	END Q[26]

	PIN Q[27]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 116.940 0.000 117.340 0.430 ;
			LAYER M1 ;
			RECT 116.940 0.000 117.340 0.430 ;
			LAYER M3 ;
			RECT 116.940 0.000 117.340 0.430 ;
		END
	END Q[27]

	PIN Q[28]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 120.830 0.000 121.230 0.430 ;
			LAYER M2 ;
			RECT 120.830 0.000 121.230 0.430 ;
			LAYER M1 ;
			RECT 120.830 0.000 121.230 0.430 ;
		END
	END Q[28]

	PIN Q[29]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 125.710 0.000 126.110 0.430 ;
			LAYER M3 ;
			RECT 125.710 0.000 126.110 0.430 ;
			LAYER M1 ;
			RECT 125.710 0.000 126.110 0.430 ;
		END
	END Q[29]

	PIN Q[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 11.940 0.000 12.340 0.430 ;
			LAYER M3 ;
			RECT 11.940 0.000 12.340 0.430 ;
			LAYER M2 ;
			RECT 11.940 0.000 12.340 0.430 ;
		END
	END Q[2]

	PIN Q[30]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 129.220 0.000 129.620 0.430 ;
			LAYER M1 ;
			RECT 129.220 0.000 129.620 0.430 ;
			LAYER M2 ;
			RECT 129.220 0.000 129.620 0.430 ;
		END
	END Q[30]

	PIN Q[31]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 133.860 0.000 134.260 0.430 ;
			LAYER M3 ;
			RECT 133.860 0.000 134.260 0.430 ;
			LAYER M1 ;
			RECT 133.860 0.000 134.260 0.430 ;
		END
	END Q[31]

	PIN Q[32]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 172.845 0.000 173.245 0.430 ;
			LAYER M3 ;
			RECT 172.845 0.000 173.245 0.430 ;
			LAYER M2 ;
			RECT 172.845 0.000 173.245 0.430 ;
		END
	END Q[32]

	PIN Q[33]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 177.095 0.000 177.495 0.430 ;
			LAYER M3 ;
			RECT 177.095 0.000 177.495 0.430 ;
			LAYER M2 ;
			RECT 177.095 0.000 177.495 0.430 ;
		END
	END Q[33]

	PIN Q[34]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 181.425 0.000 181.825 0.430 ;
			LAYER M2 ;
			RECT 181.425 0.000 181.825 0.430 ;
			LAYER M1 ;
			RECT 181.425 0.000 181.825 0.430 ;
		END
	END Q[34]

	PIN Q[35]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 185.225 0.000 185.625 0.430 ;
			LAYER M3 ;
			RECT 185.225 0.000 185.625 0.430 ;
			LAYER M1 ;
			RECT 185.225 0.000 185.625 0.430 ;
		END
	END Q[35]

	PIN Q[36]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 189.540 0.000 189.940 0.430 ;
			LAYER M2 ;
			RECT 189.540 0.000 189.940 0.430 ;
			LAYER M1 ;
			RECT 189.540 0.000 189.940 0.430 ;
		END
	END Q[36]

	PIN Q[37]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 193.740 0.000 194.140 0.430 ;
			LAYER M3 ;
			RECT 193.740 0.000 194.140 0.430 ;
			LAYER M2 ;
			RECT 193.740 0.000 194.140 0.430 ;
		END
	END Q[37]

	PIN Q[38]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 197.940 0.000 198.340 0.430 ;
			LAYER M3 ;
			RECT 197.940 0.000 198.340 0.430 ;
			LAYER M2 ;
			RECT 197.940 0.000 198.340 0.430 ;
		END
	END Q[38]

	PIN Q[39]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 202.140 0.000 202.540 0.430 ;
			LAYER M3 ;
			RECT 202.140 0.000 202.540 0.430 ;
			LAYER M2 ;
			RECT 202.140 0.000 202.540 0.430 ;
		END
	END Q[39]

	PIN Q[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 16.140 0.000 16.540 0.430 ;
			LAYER M1 ;
			RECT 16.140 0.000 16.540 0.430 ;
			LAYER M3 ;
			RECT 16.140 0.000 16.540 0.430 ;
		END
	END Q[3]

	PIN Q[40]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 206.340 0.000 206.740 0.430 ;
			LAYER M3 ;
			RECT 206.340 0.000 206.740 0.430 ;
			LAYER M2 ;
			RECT 206.340 0.000 206.740 0.430 ;
		END
	END Q[40]

	PIN Q[41]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 210.540 0.000 210.940 0.430 ;
			LAYER M3 ;
			RECT 210.540 0.000 210.940 0.430 ;
			LAYER M2 ;
			RECT 210.540 0.000 210.940 0.430 ;
		END
	END Q[41]

	PIN Q[42]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 214.740 0.000 215.140 0.430 ;
			LAYER M3 ;
			RECT 214.740 0.000 215.140 0.430 ;
			LAYER M2 ;
			RECT 214.740 0.000 215.140 0.430 ;
		END
	END Q[42]

	PIN Q[43]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 218.940 0.000 219.340 0.430 ;
			LAYER M3 ;
			RECT 218.940 0.000 219.340 0.430 ;
			LAYER M2 ;
			RECT 218.940 0.000 219.340 0.430 ;
		END
	END Q[43]

	PIN Q[44]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 223.140 0.000 223.540 0.430 ;
			LAYER M3 ;
			RECT 223.140 0.000 223.540 0.430 ;
			LAYER M2 ;
			RECT 223.140 0.000 223.540 0.430 ;
		END
	END Q[44]

	PIN Q[45]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 227.340 0.000 227.740 0.430 ;
			LAYER M3 ;
			RECT 227.340 0.000 227.740 0.430 ;
			LAYER M2 ;
			RECT 227.340 0.000 227.740 0.430 ;
		END
	END Q[45]

	PIN Q[46]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 231.540 0.000 231.940 0.430 ;
			LAYER M3 ;
			RECT 231.540 0.000 231.940 0.430 ;
			LAYER M2 ;
			RECT 231.540 0.000 231.940 0.430 ;
		END
	END Q[46]

	PIN Q[47]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 235.740 0.000 236.140 0.430 ;
			LAYER M3 ;
			RECT 235.740 0.000 236.140 0.430 ;
			LAYER M2 ;
			RECT 235.740 0.000 236.140 0.430 ;
		END
	END Q[47]

	PIN Q[48]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 239.940 0.000 240.340 0.430 ;
			LAYER M3 ;
			RECT 239.940 0.000 240.340 0.430 ;
			LAYER M2 ;
			RECT 239.940 0.000 240.340 0.430 ;
		END
	END Q[48]

	PIN Q[49]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 244.140 0.000 244.540 0.430 ;
			LAYER M2 ;
			RECT 244.140 0.000 244.540 0.430 ;
			LAYER M3 ;
			RECT 244.140 0.000 244.540 0.430 ;
		END
	END Q[49]

	PIN Q[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 20.340 0.000 20.740 0.430 ;
			LAYER M1 ;
			RECT 20.340 0.000 20.740 0.430 ;
			LAYER M3 ;
			RECT 20.340 0.000 20.740 0.430 ;
		END
	END Q[4]

	PIN Q[50]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 248.340 0.000 248.740 0.430 ;
			LAYER M2 ;
			RECT 248.340 0.000 248.740 0.430 ;
			LAYER M1 ;
			RECT 248.340 0.000 248.740 0.430 ;
		END
	END Q[50]

	PIN Q[51]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 252.540 0.000 252.940 0.430 ;
			LAYER M3 ;
			RECT 252.540 0.000 252.940 0.430 ;
			LAYER M2 ;
			RECT 252.540 0.000 252.940 0.430 ;
		END
	END Q[51]

	PIN Q[52]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 256.740 0.000 257.140 0.430 ;
			LAYER M3 ;
			RECT 256.740 0.000 257.140 0.430 ;
			LAYER M2 ;
			RECT 256.740 0.000 257.140 0.430 ;
		END
	END Q[52]

	PIN Q[53]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 260.940 0.000 261.340 0.430 ;
			LAYER M3 ;
			RECT 260.940 0.000 261.340 0.430 ;
			LAYER M2 ;
			RECT 260.940 0.000 261.340 0.430 ;
		END
	END Q[53]

	PIN Q[54]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 265.140 0.000 265.540 0.430 ;
			LAYER M3 ;
			RECT 265.140 0.000 265.540 0.430 ;
			LAYER M2 ;
			RECT 265.140 0.000 265.540 0.430 ;
		END
	END Q[54]

	PIN Q[55]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 269.340 0.000 269.740 0.430 ;
			LAYER M3 ;
			RECT 269.340 0.000 269.740 0.430 ;
			LAYER M2 ;
			RECT 269.340 0.000 269.740 0.430 ;
		END
	END Q[55]

	PIN Q[56]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 273.540 0.000 273.940 0.430 ;
			LAYER M2 ;
			RECT 273.540 0.000 273.940 0.430 ;
			LAYER M1 ;
			RECT 273.540 0.000 273.940 0.430 ;
		END
	END Q[56]

	PIN Q[57]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 277.740 0.000 278.140 0.430 ;
			LAYER M1 ;
			RECT 277.740 0.000 278.140 0.430 ;
			LAYER M2 ;
			RECT 277.740 0.000 278.140 0.430 ;
		END
	END Q[57]

	PIN Q[58]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 281.940 0.000 282.340 0.430 ;
			LAYER M1 ;
			RECT 281.940 0.000 282.340 0.430 ;
			LAYER M3 ;
			RECT 281.940 0.000 282.340 0.430 ;
		END
	END Q[58]

	PIN Q[59]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 286.140 0.000 286.540 0.430 ;
			LAYER M3 ;
			RECT 286.140 0.000 286.540 0.430 ;
			LAYER M2 ;
			RECT 286.140 0.000 286.540 0.430 ;
		END
	END Q[59]

	PIN Q[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 24.540 0.000 24.940 0.430 ;
			LAYER M2 ;
			RECT 24.540 0.000 24.940 0.430 ;
			LAYER M3 ;
			RECT 24.540 0.000 24.940 0.430 ;
		END
	END Q[5]

	PIN Q[60]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 290.340 0.000 290.740 0.430 ;
			LAYER M2 ;
			RECT 290.340 0.000 290.740 0.430 ;
			LAYER M1 ;
			RECT 290.340 0.000 290.740 0.430 ;
		END
	END Q[60]

	PIN Q[61]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 294.540 0.000 294.940 0.430 ;
			LAYER M2 ;
			RECT 294.540 0.000 294.940 0.430 ;
			LAYER M3 ;
			RECT 294.540 0.000 294.940 0.430 ;
		END
	END Q[61]

	PIN Q[62]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 298.740 0.000 299.140 0.430 ;
			LAYER M3 ;
			RECT 298.740 0.000 299.140 0.430 ;
			LAYER M2 ;
			RECT 298.740 0.000 299.140 0.430 ;
		END
	END Q[62]

	PIN Q[63]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 302.940 0.000 303.340 0.430 ;
			LAYER M3 ;
			RECT 302.940 0.000 303.340 0.430 ;
			LAYER M2 ;
			RECT 302.940 0.000 303.340 0.430 ;
		END
	END Q[63]

	PIN Q[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 28.740 0.000 29.140 0.430 ;
			LAYER M3 ;
			RECT 28.740 0.000 29.140 0.430 ;
			LAYER M2 ;
			RECT 28.740 0.000 29.140 0.430 ;
		END
	END Q[6]

	PIN Q[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 32.940 0.000 33.340 0.430 ;
			LAYER M3 ;
			RECT 32.940 0.000 33.340 0.430 ;
			LAYER M2 ;
			RECT 32.940 0.000 33.340 0.430 ;
		END
	END Q[7]

	PIN Q[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 37.140 0.000 37.540 0.430 ;
			LAYER M1 ;
			RECT 37.140 0.000 37.540 0.430 ;
			LAYER M2 ;
			RECT 37.140 0.000 37.540 0.430 ;
		END
	END Q[8]

	PIN Q[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 41.340 0.000 41.740 0.430 ;
			LAYER M1 ;
			RECT 41.340 0.000 41.740 0.430 ;
			LAYER M3 ;
			RECT 41.340 0.000 41.740 0.430 ;
		END
	END Q[9]

	PIN RTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 183.995 0.000 184.395 0.430 ;
			LAYER M1 ;
			RECT 183.995 0.000 184.395 0.430 ;
			LAYER M2 ;
			RECT 183.995 0.000 184.395 0.430 ;
		END
	END RTSEL[0]

	PIN RTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 179.305 0.000 179.705 0.430 ;
			LAYER M1 ;
			RECT 179.305 0.000 179.705 0.430 ;
			LAYER M2 ;
			RECT 179.305 0.000 179.705 0.430 ;
		END
	END RTSEL[1]

	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M4 ;
			RECT 0.500 0.000 0.830 213.850 ;
			LAYER M4 ;
			RECT 2.570 0.000 2.980 213.850 ;
			LAYER M4 ;
			RECT 6.770 0.000 7.180 213.850 ;
			LAYER M4 ;
			RECT 10.970 0.000 11.380 213.850 ;
			LAYER M4 ;
			RECT 15.170 0.000 15.580 213.850 ;
			LAYER M4 ;
			RECT 19.370 0.000 19.780 213.850 ;
			LAYER M4 ;
			RECT 23.570 0.000 23.980 213.850 ;
			LAYER M4 ;
			RECT 27.770 0.000 28.180 213.850 ;
			LAYER M4 ;
			RECT 31.970 0.000 32.380 213.850 ;
			LAYER M4 ;
			RECT 36.170 0.000 36.580 213.850 ;
			LAYER M4 ;
			RECT 40.370 0.000 40.780 213.850 ;
			LAYER M4 ;
			RECT 44.570 0.000 44.980 213.850 ;
			LAYER M4 ;
			RECT 48.770 0.000 49.180 213.850 ;
			LAYER M4 ;
			RECT 52.970 0.000 53.380 213.850 ;
			LAYER M4 ;
			RECT 57.170 0.000 57.580 213.850 ;
			LAYER M4 ;
			RECT 61.370 0.000 61.780 213.850 ;
			LAYER M4 ;
			RECT 65.570 0.000 65.980 213.850 ;
			LAYER M4 ;
			RECT 69.770 0.000 70.180 213.850 ;
			LAYER M4 ;
			RECT 73.970 0.000 74.380 213.850 ;
			LAYER M4 ;
			RECT 78.170 0.000 78.580 213.850 ;
			LAYER M4 ;
			RECT 82.370 0.000 82.780 213.850 ;
			LAYER M4 ;
			RECT 86.570 0.000 86.980 213.850 ;
			LAYER M4 ;
			RECT 90.770 0.000 91.180 213.850 ;
			LAYER M4 ;
			RECT 94.970 0.000 95.380 213.850 ;
			LAYER M4 ;
			RECT 99.170 0.000 99.580 213.850 ;
			LAYER M4 ;
			RECT 103.370 0.000 103.780 213.850 ;
			LAYER M4 ;
			RECT 107.570 0.000 107.980 213.850 ;
			LAYER M4 ;
			RECT 111.770 0.000 112.180 213.850 ;
			LAYER M4 ;
			RECT 115.970 0.000 116.380 213.850 ;
			LAYER M4 ;
			RECT 120.170 0.000 120.580 213.850 ;
			LAYER M4 ;
			RECT 124.370 0.000 124.780 213.850 ;
			LAYER M4 ;
			RECT 128.570 0.000 128.980 213.850 ;
			LAYER M4 ;
			RECT 132.770 0.000 133.180 213.850 ;
			LAYER M4 ;
			RECT 138.520 0.000 138.930 213.850 ;
			LAYER M4 ;
			RECT 147.615 0.000 148.025 213.850 ;
			LAYER M4 ;
			RECT 148.205 0.000 148.615 213.850 ;
			LAYER M4 ;
			RECT 163.665 0.000 164.075 213.850 ;
			LAYER M4 ;
			RECT 164.615 0.000 165.025 213.850 ;
			LAYER M4 ;
			RECT 171.770 0.000 172.180 213.850 ;
			LAYER M4 ;
			RECT 175.970 0.000 176.380 213.850 ;
			LAYER M4 ;
			RECT 180.170 0.000 180.580 213.850 ;
			LAYER M4 ;
			RECT 184.370 0.000 184.780 213.850 ;
			LAYER M4 ;
			RECT 188.570 0.000 188.980 213.850 ;
			LAYER M4 ;
			RECT 192.770 0.000 193.180 213.850 ;
			LAYER M4 ;
			RECT 196.970 0.000 197.380 213.850 ;
			LAYER M4 ;
			RECT 201.170 0.000 201.580 213.850 ;
			LAYER M4 ;
			RECT 205.370 0.000 205.780 213.850 ;
			LAYER M4 ;
			RECT 209.570 0.000 209.980 213.850 ;
			LAYER M4 ;
			RECT 213.770 0.000 214.180 213.850 ;
			LAYER M4 ;
			RECT 217.970 0.000 218.380 213.850 ;
			LAYER M4 ;
			RECT 222.170 0.000 222.580 213.850 ;
			LAYER M4 ;
			RECT 226.370 0.000 226.780 213.850 ;
			LAYER M4 ;
			RECT 230.570 0.000 230.980 213.850 ;
			LAYER M4 ;
			RECT 234.770 0.000 235.180 213.850 ;
			LAYER M4 ;
			RECT 238.970 0.000 239.380 213.850 ;
			LAYER M4 ;
			RECT 243.170 0.000 243.580 213.850 ;
			LAYER M4 ;
			RECT 247.370 0.000 247.780 213.850 ;
			LAYER M4 ;
			RECT 251.570 0.000 251.980 213.850 ;
			LAYER M4 ;
			RECT 255.770 0.000 256.180 213.850 ;
			LAYER M4 ;
			RECT 259.970 0.000 260.380 213.850 ;
			LAYER M4 ;
			RECT 264.170 0.000 264.580 213.850 ;
			LAYER M4 ;
			RECT 268.370 0.000 268.780 213.850 ;
			LAYER M4 ;
			RECT 272.570 0.000 272.980 213.850 ;
			LAYER M4 ;
			RECT 276.770 0.000 277.180 213.850 ;
			LAYER M4 ;
			RECT 280.970 0.000 281.380 213.850 ;
			LAYER M4 ;
			RECT 285.170 0.000 285.580 213.850 ;
			LAYER M4 ;
			RECT 289.370 0.000 289.780 213.850 ;
			LAYER M4 ;
			RECT 293.570 0.000 293.980 213.850 ;
			LAYER M4 ;
			RECT 297.770 0.000 298.180 213.850 ;
			LAYER M4 ;
			RECT 301.970 0.000 302.380 213.850 ;
			LAYER M4 ;
			RECT 306.050 0.000 306.380 213.850 ;
			LAYER M4 ;
			RECT 166.155 0.000 166.565 213.850 ;
		END
	END VDD

	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M4 ;
			RECT 5.390 0.000 6.030 213.850 ;
			LAYER M4 ;
			RECT 9.590 0.000 10.230 213.850 ;
			LAYER M4 ;
			RECT 13.790 0.000 14.430 213.850 ;
			LAYER M4 ;
			RECT 17.990 0.000 18.630 213.850 ;
			LAYER M4 ;
			RECT 22.190 0.000 22.830 213.850 ;
			LAYER M4 ;
			RECT 26.390 0.000 27.030 213.850 ;
			LAYER M4 ;
			RECT 30.590 0.000 31.230 213.850 ;
			LAYER M4 ;
			RECT 34.790 0.000 35.430 213.850 ;
			LAYER M4 ;
			RECT 38.990 0.000 39.630 213.850 ;
			LAYER M4 ;
			RECT 43.190 0.000 43.830 213.850 ;
			LAYER M4 ;
			RECT 47.390 0.000 48.030 213.850 ;
			LAYER M4 ;
			RECT 51.590 0.000 52.230 213.850 ;
			LAYER M4 ;
			RECT 55.790 0.000 56.430 213.850 ;
			LAYER M4 ;
			RECT 59.990 0.000 60.630 213.850 ;
			LAYER M4 ;
			RECT 64.190 0.000 64.830 213.850 ;
			LAYER M4 ;
			RECT 68.390 0.000 69.030 213.850 ;
			LAYER M4 ;
			RECT 72.590 0.000 73.230 213.850 ;
			LAYER M4 ;
			RECT 76.790 0.000 77.430 213.850 ;
			LAYER M4 ;
			RECT 80.990 0.000 81.630 213.850 ;
			LAYER M4 ;
			RECT 85.190 0.000 85.830 213.850 ;
			LAYER M4 ;
			RECT 89.390 0.000 90.030 213.850 ;
			LAYER M4 ;
			RECT 93.590 0.000 94.230 213.850 ;
			LAYER M4 ;
			RECT 97.790 0.000 98.430 213.850 ;
			LAYER M4 ;
			RECT 101.990 0.000 102.630 213.850 ;
			LAYER M4 ;
			RECT 106.190 0.000 106.830 213.850 ;
			LAYER M4 ;
			RECT 110.390 0.000 111.030 213.850 ;
			LAYER M4 ;
			RECT 114.590 0.000 115.230 213.850 ;
			LAYER M4 ;
			RECT 118.790 0.000 119.430 213.850 ;
			LAYER M4 ;
			RECT 122.990 0.000 123.630 213.850 ;
			LAYER M4 ;
			RECT 127.190 0.000 127.830 213.850 ;
			LAYER M4 ;
			RECT 131.390 0.000 132.030 213.850 ;
			LAYER M4 ;
			RECT 135.590 0.000 136.230 213.850 ;
			LAYER M4 ;
			RECT 137.340 0.000 137.750 213.850 ;
			LAYER M4 ;
			RECT 139.110 0.000 139.520 213.850 ;
			LAYER M4 ;
			RECT 144.665 0.000 145.075 213.850 ;
			LAYER M4 ;
			RECT 145.845 0.000 146.255 213.850 ;
			LAYER M4 ;
			RECT 147.025 0.000 147.435 213.850 ;
			LAYER M4 ;
			RECT 149.385 0.000 149.795 213.850 ;
			LAYER M4 ;
			RECT 158.225 0.000 158.635 213.850 ;
			LAYER M4 ;
			RECT 160.125 0.000 160.535 213.850 ;
			LAYER M4 ;
			RECT 162.485 0.000 162.895 213.850 ;
			LAYER M4 ;
			RECT 165.205 0.000 165.615 213.850 ;
			LAYER M4 ;
			RECT 169.005 0.000 169.415 213.850 ;
			LAYER M4 ;
			RECT 174.590 0.000 175.230 213.850 ;
			LAYER M4 ;
			RECT 178.790 0.000 179.430 213.850 ;
			LAYER M4 ;
			RECT 182.990 0.000 183.630 213.850 ;
			LAYER M4 ;
			RECT 187.190 0.000 187.830 213.850 ;
			LAYER M4 ;
			RECT 191.390 0.000 192.030 213.850 ;
			LAYER M4 ;
			RECT 195.590 0.000 196.230 213.850 ;
			LAYER M4 ;
			RECT 199.790 0.000 200.430 213.850 ;
			LAYER M4 ;
			RECT 203.990 0.000 204.630 213.850 ;
			LAYER M4 ;
			RECT 208.190 0.000 208.830 213.850 ;
			LAYER M4 ;
			RECT 212.390 0.000 213.030 213.850 ;
			LAYER M4 ;
			RECT 216.590 0.000 217.230 213.850 ;
			LAYER M4 ;
			RECT 220.790 0.000 221.430 213.850 ;
			LAYER M4 ;
			RECT 224.990 0.000 225.630 213.850 ;
			LAYER M4 ;
			RECT 229.190 0.000 229.830 213.850 ;
			LAYER M4 ;
			RECT 233.390 0.000 234.030 213.850 ;
			LAYER M4 ;
			RECT 237.590 0.000 238.230 213.850 ;
			LAYER M4 ;
			RECT 241.790 0.000 242.430 213.850 ;
			LAYER M4 ;
			RECT 245.990 0.000 246.630 213.850 ;
			LAYER M4 ;
			RECT 250.190 0.000 250.830 213.850 ;
			LAYER M4 ;
			RECT 254.390 0.000 255.030 213.850 ;
			LAYER M4 ;
			RECT 258.590 0.000 259.230 213.850 ;
			LAYER M4 ;
			RECT 262.790 0.000 263.430 213.850 ;
			LAYER M4 ;
			RECT 266.990 0.000 267.630 213.850 ;
			LAYER M4 ;
			RECT 271.190 0.000 271.830 213.850 ;
			LAYER M4 ;
			RECT 275.390 0.000 276.030 213.850 ;
			LAYER M4 ;
			RECT 279.590 0.000 280.230 213.850 ;
			LAYER M4 ;
			RECT 283.790 0.000 284.430 213.850 ;
			LAYER M4 ;
			RECT 287.990 0.000 288.630 213.850 ;
			LAYER M4 ;
			RECT 292.190 0.000 292.830 213.850 ;
			LAYER M4 ;
			RECT 296.390 0.000 297.030 213.850 ;
			LAYER M4 ;
			RECT 300.590 0.000 301.230 213.850 ;
			LAYER M4 ;
			RECT 304.790 0.000 305.430 213.850 ;
			LAYER M4 ;
			RECT 151.285 0.000 151.695 213.850 ;
			LAYER M4 ;
			RECT 161.305 0.000 161.715 213.850 ;
			LAYER M4 ;
			RECT 168.055 0.000 168.465 213.850 ;
		END
	END VSS

	PIN WEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 165.190 0.000 165.590 0.430 ;
			LAYER M3 ;
			RECT 165.190 0.000 165.590 0.430 ;
			LAYER M1 ;
			RECT 165.190 0.000 165.590 0.430 ;
		END
	END WEB

	PIN WTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 175.295 0.000 175.695 0.430 ;
			LAYER M3 ;
			RECT 175.295 0.000 175.695 0.430 ;
			LAYER M2 ;
			RECT 175.295 0.000 175.695 0.430 ;
		END
	END WTSEL[0]

	PIN WTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 171.045 0.000 171.445 0.430 ;
			LAYER M2 ;
			RECT 171.045 0.000 171.445 0.430 ;
			LAYER M3 ;
			RECT 171.045 0.000 171.445 0.430 ;
		END
	END WTSEL[1]

	PIN WTSEL[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 173.445 0.000 173.845 0.430 ;
			LAYER M1 ;
			RECT 173.445 0.000 173.845 0.430 ;
			LAYER M2 ;
			RECT 173.445 0.000 173.845 0.430 ;
		END
	END WTSEL[2]
	OBS
		# Promoted blockages
		LAYER M3 ;
		RECT 265.690 0.000 266.190 0.430 ;
		LAYER M2 ;
		RECT 265.690 0.000 266.190 0.430 ;
		LAYER M1 ;
		RECT 274.080 0.000 274.600 0.430 ;
		LAYER M1 ;
		RECT 271.080 0.000 272.200 0.430 ;
		LAYER M2 ;
		RECT 269.890 0.000 270.390 0.430 ;
		LAYER M1 ;
		RECT 298.080 0.000 298.600 0.430 ;
		LAYER VIA3 ;
		RECT 298.090 0.000 298.590 0.430 ;
		LAYER M2 ;
		RECT 298.090 0.000 298.590 0.430 ;
		LAYER VIA3 ;
		RECT 296.290 0.000 297.390 0.430 ;
		LAYER M3 ;
		RECT 296.290 0.000 297.390 0.430 ;
		LAYER M3 ;
		RECT 298.090 0.000 298.590 0.430 ;
		LAYER M1 ;
		RECT 299.280 0.000 299.800 0.430 ;
		LAYER M2 ;
		RECT 286.690 0.000 287.190 0.430 ;
		LAYER M2 ;
		RECT 287.890 0.000 288.990 0.430 ;
		LAYER M1 ;
		RECT 292.080 0.000 293.200 0.430 ;
		LAYER M1 ;
		RECT 296.280 0.000 297.400 0.430 ;
		LAYER VIA3 ;
		RECT 299.290 0.000 299.790 0.430 ;
		LAYER M1 ;
		RECT 264.480 0.000 265.000 0.430 ;
		LAYER VIA3 ;
		RECT 264.490 0.000 264.990 0.430 ;
		LAYER VIA3 ;
		RECT 265.690 0.000 266.190 0.430 ;
		LAYER VIA3 ;
		RECT 269.890 0.000 270.390 0.430 ;
		LAYER M1 ;
		RECT 269.880 0.000 270.400 0.430 ;
		LAYER M2 ;
		RECT 285.490 0.000 285.990 0.430 ;
		LAYER M1 ;
		RECT 285.480 0.000 286.000 0.430 ;
		LAYER M1 ;
		RECT 286.680 0.000 287.200 0.430 ;
		LAYER M2 ;
		RECT 283.690 0.000 284.790 0.430 ;
		LAYER VIA3 ;
		RECT 290.890 0.000 291.390 0.430 ;
		LAYER M2 ;
		RECT 290.890 0.000 291.390 0.430 ;
		LAYER M2 ;
		RECT 289.690 0.000 290.190 0.430 ;
		LAYER M3 ;
		RECT 289.690 0.000 290.190 0.430 ;
		LAYER M3 ;
		RECT 287.890 0.000 288.990 0.430 ;
		LAYER M1 ;
		RECT 287.880 0.000 289.000 0.430 ;
		LAYER VIA3 ;
		RECT 295.090 0.000 295.590 0.430 ;
		LAYER M3 ;
		RECT 295.090 0.000 295.590 0.430 ;
		LAYER VIA3 ;
		RECT 293.890 0.000 294.390 0.430 ;
		LAYER M2 ;
		RECT 295.090 0.000 295.590 0.430 ;
		LAYER M2 ;
		RECT 281.290 0.000 281.790 0.430 ;
		LAYER M2 ;
		RECT 282.490 0.000 282.990 0.430 ;
		LAYER VIA3 ;
		RECT 277.090 0.000 277.590 0.430 ;
		LAYER M3 ;
		RECT 285.490 0.000 285.990 0.430 ;
		LAYER VIA3 ;
		RECT 285.490 0.000 285.990 0.430 ;
		LAYER M1 ;
		RECT 283.680 0.000 284.800 0.430 ;
		LAYER M2 ;
		RECT 300.490 0.000 301.590 0.430 ;
		LAYER M1 ;
		RECT 300.480 0.000 301.600 0.430 ;
		LAYER M2 ;
		RECT 302.290 0.000 302.790 0.430 ;
		LAYER M3 ;
		RECT 302.290 0.000 302.790 0.430 ;
		LAYER VIA3 ;
		RECT 300.490 0.000 301.590 0.430 ;
		LAYER M3 ;
		RECT 300.490 0.000 301.590 0.430 ;
		LAYER M1 ;
		RECT 302.280 0.000 302.800 0.430 ;
		LAYER VIA3 ;
		RECT 302.290 0.000 302.790 0.430 ;
		LAYER M3 ;
		RECT 303.490 0.000 303.990 0.430 ;
		LAYER VIA3 ;
		RECT 303.490 0.000 303.990 0.430 ;
		LAYER M2 ;
		RECT 296.290 0.000 297.390 0.430 ;
		LAYER M3 ;
		RECT 293.890 0.000 294.390 0.430 ;
		LAYER M1 ;
		RECT 295.080 0.000 295.600 0.430 ;
		LAYER M2 ;
		RECT 293.890 0.000 294.390 0.430 ;
		LAYER M1 ;
		RECT 290.880 0.000 291.400 0.430 ;
		LAYER M3 ;
		RECT 290.890 0.000 291.390 0.430 ;
		LAYER M2 ;
		RECT 292.090 0.000 293.190 0.430 ;
		LAYER M3 ;
		RECT 292.090 0.000 293.190 0.430 ;
		LAYER VIA3 ;
		RECT 292.090 0.000 293.190 0.430 ;
		LAYER M4 ;
		RECT 281.380 0.000 283.790 213.850 ;
		LAYER M4 ;
		RECT 267.630 0.000 268.370 213.850 ;
		LAYER M4 ;
		RECT 271.830 0.000 272.570 213.850 ;
		LAYER M4 ;
		RECT 268.780 0.000 271.190 213.850 ;
		LAYER M4 ;
		RECT 293.980 0.000 296.390 213.850 ;
		LAYER M4 ;
		RECT 292.830 0.000 293.570 213.850 ;
		LAYER M4 ;
		RECT 285.580 0.000 287.990 213.850 ;
		LAYER M4 ;
		RECT 284.430 0.000 285.170 213.850 ;
		LAYER M4 ;
		RECT 289.780 0.000 292.190 213.850 ;
		LAYER M4 ;
		RECT 288.630 0.000 289.370 213.850 ;
		LAYER M4 ;
		RECT 302.380 0.000 304.790 213.850 ;
		LAYER M4 ;
		RECT 301.230 0.000 301.970 213.850 ;
		LAYER M4 ;
		RECT 298.180 0.000 300.590 213.850 ;
		LAYER M4 ;
		RECT 297.030 0.000 297.770 213.850 ;
		LAYER M4 ;
		RECT 305.430 0.000 306.050 213.850 ;
		LAYER M4 ;
		RECT 264.580 0.000 266.990 213.850 ;
		LAYER M4 ;
		RECT 263.430 0.000 264.170 213.850 ;
		LAYER M4 ;
		RECT 280.230 0.000 280.970 213.850 ;
		LAYER M4 ;
		RECT 277.180 0.000 279.590 213.850 ;
		LAYER M4 ;
		RECT 276.030 0.000 276.770 213.850 ;
		LAYER M4 ;
		RECT 272.980 0.000 275.390 213.850 ;
		LAYER M1 ;
		RECT 281.280 0.000 281.800 0.430 ;
		LAYER M3 ;
		RECT 281.290 0.000 281.790 0.430 ;
		LAYER VIA3 ;
		RECT 283.690 0.000 284.790 0.430 ;
		LAYER M2 ;
		RECT 279.490 0.000 280.590 0.430 ;
		LAYER M3 ;
		RECT 304.690 0.000 306.880 0.430 ;
		LAYER VIA3 ;
		RECT 304.690 0.000 306.880 0.430 ;
		LAYER M1 ;
		RECT 303.480 0.000 304.000 0.430 ;
		LAYER VIA3 ;
		RECT 281.290 0.000 281.790 0.430 ;
		LAYER M1 ;
		RECT 293.880 0.000 294.400 0.430 ;
		LAYER VIA3 ;
		RECT 287.890 0.000 288.990 0.430 ;
		LAYER M1 ;
		RECT 289.680 0.000 290.200 0.430 ;
		LAYER VIA3 ;
		RECT 289.690 0.000 290.190 0.430 ;
		LAYER M3 ;
		RECT 282.490 0.000 282.990 0.430 ;
		LAYER VIA3 ;
		RECT 282.490 0.000 282.990 0.430 ;
		LAYER M1 ;
		RECT 282.480 0.000 283.000 0.430 ;
		LAYER M3 ;
		RECT 283.690 0.000 284.790 0.430 ;
		LAYER M4 ;
		RECT 256.180 0.000 258.590 213.850 ;
		LAYER M4 ;
		RECT 255.030 0.000 255.770 213.850 ;
		LAYER M4 ;
		RECT 251.980 0.000 254.390 213.850 ;
		LAYER M4 ;
		RECT 250.830 0.000 251.570 213.850 ;
		LAYER VIA3 ;
		RECT 220.690 0.000 221.790 0.430 ;
		LAYER M3 ;
		RECT 216.490 0.000 217.590 0.430 ;
		LAYER M2 ;
		RECT 216.490 0.000 217.590 0.430 ;
		LAYER M4 ;
		RECT 225.630 0.000 226.370 213.850 ;
		LAYER M4 ;
		RECT 247.780 0.000 250.190 213.850 ;
		LAYER M4 ;
		RECT 246.630 0.000 247.370 213.850 ;
		LAYER M4 ;
		RECT 243.580 0.000 245.990 213.850 ;
		LAYER M4 ;
		RECT 242.430 0.000 243.170 213.850 ;
		LAYER M4 ;
		RECT 239.380 0.000 241.790 213.850 ;
		LAYER M2 ;
		RECT 218.290 0.000 218.790 0.430 ;
		LAYER M3 ;
		RECT 218.290 0.000 218.790 0.430 ;
		LAYER VIA3 ;
		RECT 219.490 0.000 219.990 0.430 ;
		LAYER M3 ;
		RECT 219.490 0.000 219.990 0.430 ;
		LAYER VIA3 ;
		RECT 215.290 0.000 215.790 0.430 ;
		LAYER M1 ;
		RECT 214.080 0.000 214.600 0.430 ;
		LAYER M2 ;
		RECT 212.290 0.000 213.390 0.430 ;
		LAYER VIA3 ;
		RECT 211.090 0.000 211.590 0.430 ;
		LAYER M3 ;
		RECT 209.890 0.000 210.390 0.430 ;
		LAYER VIA3 ;
		RECT 209.890 0.000 210.390 0.430 ;
		LAYER M1 ;
		RECT 216.480 0.000 217.600 0.430 ;
		LAYER M4 ;
		RECT 213.030 0.000 213.770 213.850 ;
		LAYER M3 ;
		RECT 211.090 0.000 211.590 0.430 ;
		LAYER M4 ;
		RECT 209.980 0.000 212.390 213.850 ;
		LAYER M4 ;
		RECT 201.580 0.000 203.990 213.850 ;
		LAYER M1 ;
		RECT 304.680 0.000 306.880 0.430 ;
		LAYER M2 ;
		RECT 303.490 0.000 303.990 0.430 ;
		LAYER M2 ;
		RECT 299.290 0.000 299.790 0.430 ;
		LAYER M3 ;
		RECT 299.290 0.000 299.790 0.430 ;
		LAYER M2 ;
		RECT 16.690 0.000 17.190 0.430 ;
		LAYER M3 ;
		RECT 16.690 0.000 17.190 0.430 ;
		LAYER VIA3 ;
		RECT 16.690 0.000 17.190 0.430 ;
		LAYER M1 ;
		RECT 16.680 0.000 17.200 0.430 ;
		LAYER M2 ;
		RECT 15.490 0.000 15.990 0.430 ;
		LAYER M1 ;
		RECT 15.480 0.000 16.000 0.430 ;
		LAYER M2 ;
		RECT 211.090 0.000 211.590 0.430 ;
		LAYER M4 ;
		RECT 0.830 0.000 1.450 213.850 ;
		LAYER M4 ;
		RECT 1.830 0.000 2.570 213.850 ;
		LAYER M2 ;
		RECT 0.000 0.000 2.190 213.850 ;
		LAYER M3 ;
		RECT 0.000 0.000 2.190 213.850 ;
		LAYER VIA3 ;
		RECT 0.000 0.000 2.190 213.850 ;
		LAYER M1 ;
		RECT 0.000 0.000 2.200 213.850 ;
		LAYER M4 ;
		RECT 200.430 0.000 201.170 213.850 ;
		LAYER VIA3 ;
		RECT 2.190 0.430 306.880 213.850 ;
		LAYER M2 ;
		RECT 2.190 0.430 306.880 213.850 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 306.880 213.850 ;
		LAYER M4 ;
		RECT 7.180 0.000 9.590 213.850 ;
		LAYER M3 ;
		RECT 2.190 0.430 306.880 213.850 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 306.880 213.850 ;
		LAYER M4 ;
		RECT 15.580 0.000 17.990 213.850 ;
		LAYER M4 ;
		RECT 14.430 0.000 15.170 213.850 ;
		LAYER M4 ;
		RECT 11.380 0.000 13.790 213.850 ;
		LAYER M4 ;
		RECT 10.230 0.000 10.970 213.850 ;
		LAYER M4 ;
		RECT 2.980 0.000 5.390 213.850 ;
		LAYER M4 ;
		RECT 6.030 0.000 6.770 213.850 ;
		LAYER M1 ;
		RECT 2.200 0.430 306.880 213.850 ;
		LAYER M4 ;
		RECT 196.230 0.000 196.970 213.850 ;
		LAYER M5 ;
		RECT 0.000 0.000 306.880 0.100 ;
		LAYER M5 ;
		RECT 0.000 213.750 306.880 213.850 ;
		LAYER M4 ;
		RECT 187.830 0.000 188.570 213.850 ;
		LAYER M4 ;
		RECT 184.780 0.000 187.190 213.850 ;
		LAYER M4 ;
		RECT 183.630 0.000 184.370 213.850 ;
		LAYER M4 ;
		RECT 136.340 0.000 137.340 213.850 ;
		LAYER M4 ;
		RECT 115.230 0.000 115.970 213.850 ;
		LAYER M4 ;
		RECT 112.180 0.000 114.590 213.850 ;
		LAYER M4 ;
		RECT 111.030 0.000 111.770 213.850 ;
		LAYER M4 ;
		RECT 138.930 0.000 139.110 213.850 ;
		LAYER M4 ;
		RECT 137.750 0.000 138.520 213.850 ;
		LAYER M4 ;
		RECT 132.030 0.000 132.770 213.850 ;
		LAYER M4 ;
		RECT 128.980 0.000 131.390 213.850 ;
		LAYER M4 ;
		RECT 127.830 0.000 128.570 213.850 ;
		LAYER M4 ;
		RECT 124.780 0.000 127.190 213.850 ;
		LAYER M4 ;
		RECT 133.180 0.000 135.590 213.850 ;
		LAYER M4 ;
		RECT 116.380 0.000 118.790 213.850 ;
		LAYER M4 ;
		RECT 120.580 0.000 122.990 213.850 ;
		LAYER M4 ;
		RECT 123.630 0.000 124.370 213.850 ;
		LAYER M4 ;
		RECT 119.430 0.000 120.170 213.850 ;
		LAYER M4 ;
		RECT 149.795 0.000 151.285 213.850 ;
		LAYER M4 ;
		RECT 146.255 0.000 147.025 213.850 ;
		LAYER M4 ;
		RECT 145.075 0.000 145.845 213.850 ;
		LAYER M4 ;
		RECT 139.520 0.000 144.665 213.850 ;
		LAYER M4 ;
		RECT 188.980 0.000 191.390 213.850 ;
		LAYER M4 ;
		RECT 192.030 0.000 192.770 213.850 ;
		LAYER M4 ;
		RECT 193.180 0.000 195.590 213.850 ;
		LAYER M4 ;
		RECT 197.380 0.000 199.790 213.850 ;
		LAYER M4 ;
		RECT 107.980 0.000 110.390 213.850 ;
		LAYER M4 ;
		RECT 91.180 0.000 93.590 213.850 ;
		LAYER M4 ;
		RECT 90.030 0.000 90.770 213.850 ;
		LAYER M4 ;
		RECT 74.380 0.000 76.790 213.850 ;
		LAYER M4 ;
		RECT 106.830 0.000 107.570 213.850 ;
		LAYER M4 ;
		RECT 102.630 0.000 103.370 213.850 ;
		LAYER M4 ;
		RECT 95.380 0.000 97.790 213.850 ;
		LAYER M4 ;
		RECT 94.230 0.000 94.970 213.850 ;
		LAYER M4 ;
		RECT 260.380 0.000 262.790 213.850 ;
		LAYER M4 ;
		RECT 69.030 0.000 69.770 213.850 ;
		LAYER M4 ;
		RECT 35.430 0.000 36.170 213.850 ;
		LAYER M4 ;
		RECT 73.230 0.000 73.970 213.850 ;
		LAYER M1 ;
		RECT 208.080 0.000 209.200 0.430 ;
		LAYER M2 ;
		RECT 57.490 0.000 57.990 0.430 ;
		LAYER M3 ;
		RECT 57.490 0.000 57.990 0.430 ;
		LAYER M3 ;
		RECT 58.690 0.000 59.190 0.430 ;
		LAYER VIA3 ;
		RECT 58.690 0.000 59.190 0.430 ;
		LAYER M2 ;
		RECT 58.690 0.000 59.190 0.430 ;
		LAYER M3 ;
		RECT 59.890 0.000 60.990 0.430 ;
		LAYER M2 ;
		RECT 49.090 0.000 49.590 0.430 ;
		LAYER M2 ;
		RECT 55.690 0.000 56.790 0.430 ;
		LAYER M1 ;
		RECT 54.480 0.000 55.000 0.430 ;
		LAYER M3 ;
		RECT 36.490 0.000 36.990 0.430 ;
		LAYER M2 ;
		RECT 37.690 0.000 38.190 0.430 ;
		LAYER M3 ;
		RECT 37.690 0.000 38.190 0.430 ;
		LAYER M3 ;
		RECT 198.490 0.000 198.990 0.430 ;
		LAYER M2 ;
		RECT 68.290 0.000 69.390 0.430 ;
		LAYER M3 ;
		RECT 64.090 0.000 65.190 0.430 ;
		LAYER M1 ;
		RECT 93.480 0.000 94.600 0.430 ;
		LAYER M3 ;
		RECT 92.290 0.000 92.790 0.430 ;
		LAYER VIA3 ;
		RECT 92.290 0.000 92.790 0.430 ;
		LAYER M1 ;
		RECT 32.280 0.000 32.800 0.430 ;
		LAYER M2 ;
		RECT 32.290 0.000 32.790 0.430 ;
		LAYER M3 ;
		RECT 32.290 0.000 32.790 0.430 ;
		LAYER M1 ;
		RECT 33.480 0.000 34.000 0.430 ;
		LAYER M3 ;
		RECT 33.490 0.000 33.990 0.430 ;
		LAYER M2 ;
		RECT 33.490 0.000 33.990 0.430 ;
		LAYER M2 ;
		RECT 34.690 0.000 35.790 0.430 ;
		LAYER M1 ;
		RECT 34.680 0.000 35.800 0.430 ;
		LAYER VIA3 ;
		RECT 33.490 0.000 33.990 0.430 ;
		LAYER M2 ;
		RECT 38.890 0.000 39.990 0.430 ;
		LAYER M1 ;
		RECT 38.880 0.000 40.000 0.430 ;
		LAYER VIA3 ;
		RECT 41.890 0.000 42.390 0.430 ;
		LAYER M2 ;
		RECT 43.090 0.000 44.190 0.430 ;
		LAYER M3 ;
		RECT 43.090 0.000 44.190 0.430 ;
		LAYER VIA3 ;
		RECT 37.690 0.000 38.190 0.430 ;
		LAYER M2 ;
		RECT 36.490 0.000 36.990 0.430 ;
		LAYER VIA3 ;
		RECT 36.490 0.000 36.990 0.430 ;
		LAYER M4 ;
		RECT 180.580 0.000 182.990 213.850 ;
		LAYER M4 ;
		RECT 179.430 0.000 180.170 213.850 ;
		LAYER M4 ;
		RECT 176.380 0.000 178.790 213.850 ;
		LAYER M4 ;
		RECT 175.230 0.000 175.970 213.850 ;
		LAYER M4 ;
		RECT 169.415 30.270 171.030 120.760 ;
		LAYER M4 ;
		RECT 171.030 27.670 171.770 120.760 ;
		LAYER M4 ;
		RECT 172.180 0.000 174.590 213.850 ;
		LAYER M4 ;
		RECT 169.415 120.760 171.770 213.850 ;
		LAYER M4 ;
		RECT 169.415 0.000 171.770 30.270 ;
		LAYER M4 ;
		RECT 168.465 0.000 169.005 213.850 ;
		LAYER M4 ;
		RECT 166.565 0.000 168.055 213.850 ;
		LAYER M4 ;
		RECT 165.615 0.000 166.155 213.850 ;
		LAYER M4 ;
		RECT 148.615 0.000 149.385 213.850 ;
		LAYER M4 ;
		RECT 148.025 0.000 148.205 213.850 ;
		LAYER M4 ;
		RECT 147.435 0.000 147.615 213.850 ;
		LAYER M4 ;
		RECT 158.635 0.000 160.125 213.850 ;
		LAYER M4 ;
		RECT 165.025 0.000 165.205 213.850 ;
		LAYER M4 ;
		RECT 151.695 0.000 158.225 213.850 ;
		LAYER M4 ;
		RECT 160.535 0.000 161.305 213.850 ;
		LAYER M4 ;
		RECT 161.715 0.000 162.485 213.850 ;
		LAYER M4 ;
		RECT 162.895 0.000 163.665 213.850 ;
		LAYER M4 ;
		RECT 164.075 0.000 164.615 213.850 ;
		LAYER M4 ;
		RECT 205.780 0.000 208.190 213.850 ;
		LAYER M4 ;
		RECT 229.830 0.000 230.570 213.850 ;
		LAYER M4 ;
		RECT 221.430 0.000 222.170 213.850 ;
		LAYER M4 ;
		RECT 226.780 0.000 229.190 213.850 ;
		LAYER M4 ;
		RECT 222.580 0.000 224.990 213.850 ;
		LAYER M4 ;
		RECT 208.830 0.000 209.570 213.850 ;
		LAYER M4 ;
		RECT 214.180 0.000 216.590 213.850 ;
		LAYER M4 ;
		RECT 217.230 0.000 217.970 213.850 ;
		LAYER M4 ;
		RECT 218.380 0.000 220.790 213.850 ;
		LAYER M4 ;
		RECT 204.630 0.000 205.370 213.850 ;
		LAYER M4 ;
		RECT 234.030 0.000 234.770 213.850 ;
		LAYER M4 ;
		RECT 230.980 0.000 233.390 213.850 ;
		LAYER M4 ;
		RECT 259.230 0.000 259.970 213.850 ;
		LAYER M4 ;
		RECT 235.180 0.000 237.590 213.850 ;
		LAYER M4 ;
		RECT 238.230 0.000 238.970 213.850 ;
		LAYER M4 ;
		RECT 61.780 0.000 64.190 213.850 ;
		LAYER M4 ;
		RECT 64.830 0.000 65.570 213.850 ;
		LAYER M4 ;
		RECT 65.980 0.000 68.390 213.850 ;
		LAYER M4 ;
		RECT 70.180 0.000 72.590 213.850 ;
		LAYER M4 ;
		RECT 60.630 0.000 61.370 213.850 ;
		LAYER M4 ;
		RECT 52.230 0.000 52.970 213.850 ;
		LAYER M4 ;
		RECT 53.380 0.000 55.790 213.850 ;
		LAYER M4 ;
		RECT 56.430 0.000 57.170 213.850 ;
		LAYER M4 ;
		RECT 57.580 0.000 59.990 213.850 ;
		LAYER M4 ;
		RECT 48.030 0.000 48.770 213.850 ;
		LAYER M4 ;
		RECT 49.180 0.000 51.590 213.850 ;
		LAYER M4 ;
		RECT 77.430 0.000 78.170 213.850 ;
		LAYER M4 ;
		RECT 40.780 0.000 43.190 213.850 ;
		LAYER M4 ;
		RECT 43.830 0.000 44.570 213.850 ;
		LAYER M4 ;
		RECT 44.980 0.000 47.390 213.850 ;
		LAYER M4 ;
		RECT 86.980 0.000 89.390 213.850 ;
		LAYER M4 ;
		RECT 98.430 0.000 99.170 213.850 ;
		LAYER M4 ;
		RECT 99.580 0.000 101.990 213.850 ;
		LAYER M4 ;
		RECT 103.780 0.000 106.190 213.850 ;
		LAYER M4 ;
		RECT 85.830 0.000 86.570 213.850 ;
		LAYER M4 ;
		RECT 82.780 0.000 85.190 213.850 ;
		LAYER M4 ;
		RECT 81.630 0.000 82.370 213.850 ;
		LAYER M4 ;
		RECT 78.580 0.000 80.990 213.850 ;
		LAYER M4 ;
		RECT 39.630 0.000 40.370 213.850 ;
		LAYER M4 ;
		RECT 36.580 0.000 38.990 213.850 ;
		LAYER M4 ;
		RECT 18.630 0.000 19.370 213.850 ;
		LAYER M4 ;
		RECT 32.380 0.000 34.790 213.850 ;
		LAYER M4 ;
		RECT 31.230 0.000 31.970 213.850 ;
		LAYER M4 ;
		RECT 19.780 0.000 22.190 213.850 ;
		LAYER M4 ;
		RECT 28.180 0.000 30.590 213.850 ;
		LAYER M4 ;
		RECT 27.030 0.000 27.770 213.850 ;
		LAYER M4 ;
		RECT 23.980 0.000 26.390 213.850 ;
		LAYER M4 ;
		RECT 22.830 0.000 23.570 213.850 ;
		LAYER M2 ;
		RECT 304.690 0.000 306.880 0.430 ;
		LAYER M3 ;
		RECT 286.690 0.000 287.190 0.430 ;
		LAYER VIA3 ;
		RECT 286.690 0.000 287.190 0.430 ;
		LAYER M2 ;
		RECT 219.490 0.000 219.990 0.430 ;
		LAYER VIA3 ;
		RECT 218.290 0.000 218.790 0.430 ;
		LAYER M1 ;
		RECT 218.280 0.000 218.800 0.430 ;
		LAYER VIA3 ;
		RECT 214.090 0.000 214.590 0.430 ;
		LAYER M3 ;
		RECT 220.690 0.000 221.790 0.430 ;
		LAYER M3 ;
		RECT 212.290 0.000 213.390 0.430 ;
		LAYER M1 ;
		RECT 212.280 0.000 213.400 0.430 ;
		LAYER M2 ;
		RECT 209.890 0.000 210.390 0.430 ;
		LAYER M2 ;
		RECT 17.890 0.000 18.990 0.430 ;
		LAYER M3 ;
		RECT 17.890 0.000 18.990 0.430 ;
		LAYER M1 ;
		RECT 30.480 0.000 31.600 0.430 ;
		LAYER M3 ;
		RECT 30.490 0.000 31.590 0.430 ;
		LAYER VIA3 ;
		RECT 30.490 0.000 31.590 0.430 ;
		LAYER M2 ;
		RECT 19.690 0.000 20.190 0.430 ;
		LAYER M2 ;
		RECT 29.290 0.000 29.790 0.430 ;
		LAYER M2 ;
		RECT 20.890 0.000 21.390 0.430 ;
		LAYER M1 ;
		RECT 118.680 0.000 119.490 0.430 ;
		LAYER M3 ;
		RECT 117.490 0.000 117.990 0.430 ;
		LAYER VIA3 ;
		RECT 117.490 0.000 117.990 0.430 ;
		LAYER M2 ;
		RECT 117.490 0.000 117.990 0.430 ;
		LAYER VIA3 ;
		RECT 118.690 0.000 119.480 0.430 ;
		LAYER M2 ;
		RECT 120.180 0.000 120.680 0.430 ;
		LAYER M3 ;
		RECT 120.180 0.000 120.680 0.430 ;
		LAYER M1 ;
		RECT 120.170 0.000 120.690 0.430 ;
		LAYER M1 ;
		RECT 121.370 0.000 122.570 0.430 ;
		LAYER VIA3 ;
		RECT 120.180 0.000 120.680 0.430 ;
		LAYER M3 ;
		RECT 121.380 0.000 122.560 0.430 ;
		LAYER M2 ;
		RECT 123.260 0.000 123.670 0.430 ;
		LAYER M3 ;
		RECT 123.260 0.000 123.670 0.430 ;
		LAYER VIA3 ;
		RECT 123.260 0.000 123.670 0.430 ;
		LAYER M3 ;
		RECT 118.690 0.000 119.480 0.430 ;
		LAYER M2 ;
		RECT 118.690 0.000 119.480 0.430 ;
		LAYER M1 ;
		RECT 117.480 0.000 118.000 0.430 ;
		LAYER M2 ;
		RECT 124.370 0.000 125.560 0.430 ;
		LAYER M3 ;
		RECT 124.370 0.000 125.560 0.430 ;
		LAYER VIA3 ;
		RECT 124.370 0.000 125.560 0.430 ;
		LAYER M2 ;
		RECT 121.380 0.000 122.560 0.430 ;
		LAYER VIA3 ;
		RECT 121.380 0.000 122.560 0.430 ;
		LAYER M1 ;
		RECT 123.250 0.000 123.680 0.430 ;
		LAYER M1 ;
		RECT 128.190 0.000 129.080 0.430 ;
		LAYER M3 ;
		RECT 129.770 0.000 130.520 0.430 ;
		LAYER VIA3 ;
		RECT 129.770 0.000 130.520 0.430 ;
		LAYER M1 ;
		RECT 129.760 0.000 130.530 0.430 ;
		LAYER VIA3 ;
		RECT 135.710 0.000 138.020 0.430 ;
		LAYER M3 ;
		RECT 135.710 0.000 138.020 0.430 ;
		LAYER M1 ;
		RECT 132.420 0.000 133.720 0.430 ;
		LAYER M2 ;
		RECT 135.710 0.000 138.020 0.430 ;
		LAYER M1 ;
		RECT 135.700 0.000 138.030 0.430 ;
		LAYER M3 ;
		RECT 134.410 0.000 135.010 0.430 ;
		LAYER M1 ;
		RECT 134.400 0.000 135.020 0.430 ;
		LAYER M1 ;
		RECT 142.470 0.000 142.490 0.430 ;
		LAYER M3 ;
		RECT 139.420 0.000 141.780 0.430 ;
		LAYER M2 ;
		RECT 139.420 0.000 141.780 0.430 ;
		LAYER M1 ;
		RECT 139.410 0.000 141.790 0.430 ;
		LAYER VIA3 ;
		RECT 139.420 0.000 141.780 0.430 ;
		LAYER M2 ;
		RECT 143.180 0.000 145.540 0.430 ;
		LAYER M3 ;
		RECT 131.220 0.000 131.730 0.430 ;
		LAYER M2 ;
		RECT 131.220 0.000 131.730 0.430 ;
		LAYER VIA3 ;
		RECT 131.220 0.000 131.730 0.430 ;
		LAYER M1 ;
		RECT 116.280 0.000 116.800 0.430 ;
		LAYER M3 ;
		RECT 126.260 0.000 126.830 0.430 ;
		LAYER M1 ;
		RECT 124.360 0.000 125.570 0.430 ;
		LAYER VIA3 ;
		RECT 126.260 0.000 126.830 0.430 ;
		LAYER M2 ;
		RECT 126.260 0.000 126.830 0.430 ;
		LAYER M1 ;
		RECT 126.250 0.000 126.840 0.430 ;
		LAYER M2 ;
		RECT 134.410 0.000 135.010 0.430 ;
		LAYER M3 ;
		RECT 132.430 0.000 133.710 0.430 ;
		LAYER VIA3 ;
		RECT 132.430 0.000 133.710 0.430 ;
		LAYER M2 ;
		RECT 132.430 0.000 133.710 0.430 ;
		LAYER M1 ;
		RECT 143.170 0.000 145.550 0.430 ;
		LAYER M1 ;
		RECT 146.230 0.000 146.250 0.430 ;
		LAYER M1 ;
		RECT 138.710 0.000 138.730 0.430 ;
		LAYER M1 ;
		RECT 146.930 0.000 153.070 0.430 ;
		LAYER M3 ;
		RECT 143.180 0.000 145.540 0.430 ;
		LAYER VIA3 ;
		RECT 143.180 0.000 145.540 0.430 ;
		LAYER VIA3 ;
		RECT 134.410 0.000 135.010 0.430 ;
		LAYER M1 ;
		RECT 131.210 0.000 131.740 0.430 ;
		LAYER M2 ;
		RECT 129.770 0.000 130.520 0.430 ;
		LAYER VIA3 ;
		RECT 128.200 0.000 129.070 0.430 ;
		LAYER M2 ;
		RECT 128.200 0.000 129.070 0.430 ;
		LAYER M3 ;
		RECT 128.200 0.000 129.070 0.430 ;
		LAYER M2 ;
		RECT 153.760 0.000 156.820 0.430 ;
		LAYER M1 ;
		RECT 153.750 0.000 156.830 0.430 ;
		LAYER M1 ;
		RECT 157.510 0.000 157.530 0.430 ;
		LAYER M2 ;
		RECT 146.940 0.000 153.060 0.430 ;
		LAYER M3 ;
		RECT 153.760 0.000 156.820 0.430 ;
		LAYER VIA3 ;
		RECT 153.760 0.000 156.820 0.430 ;
		LAYER M3 ;
		RECT 146.940 0.000 153.060 0.430 ;
		LAYER VIA3 ;
		RECT 146.940 0.000 153.060 0.430 ;
		LAYER M1 ;
		RECT 59.880 0.000 61.000 0.430 ;
		LAYER M1 ;
		RECT 68.280 0.000 69.400 0.430 ;
		LAYER M3 ;
		RECT 68.290 0.000 69.390 0.430 ;
		LAYER M2 ;
		RECT 61.690 0.000 62.190 0.430 ;
		LAYER VIA3 ;
		RECT 67.090 0.000 67.590 0.430 ;
		LAYER M3 ;
		RECT 67.090 0.000 67.590 0.430 ;
		LAYER M1 ;
		RECT 70.080 0.000 70.600 0.430 ;
		LAYER M2 ;
		RECT 89.290 0.000 90.390 0.430 ;
		LAYER M1 ;
		RECT 91.080 0.000 91.600 0.430 ;
		LAYER VIA3 ;
		RECT 70.090 0.000 70.590 0.430 ;
		LAYER M1 ;
		RECT 92.280 0.000 92.800 0.430 ;
		LAYER M3 ;
		RECT 93.490 0.000 94.590 0.430 ;
		LAYER M2 ;
		RECT 92.290 0.000 92.790 0.430 ;
		LAYER VIA3 ;
		RECT 93.490 0.000 94.590 0.430 ;
		LAYER M3 ;
		RECT 208.090 0.000 209.190 0.430 ;
		LAYER M1 ;
		RECT 215.280 0.000 215.800 0.430 ;
		LAYER VIA3 ;
		RECT 216.490 0.000 217.590 0.430 ;
		LAYER M1 ;
		RECT 219.480 0.000 220.000 0.430 ;
		LAYER M3 ;
		RECT 180.455 0.000 181.275 0.430 ;
		LAYER M3 ;
		RECT 173.995 0.000 174.495 0.430 ;
		LAYER VIA3 ;
		RECT 173.995 0.000 174.495 0.430 ;
		LAYER M2 ;
		RECT 173.995 0.000 174.495 0.430 ;
		LAYER M2 ;
		RECT 197.290 0.000 197.790 0.430 ;
		LAYER M1 ;
		RECT 170.120 0.000 170.905 0.430 ;
		LAYER M3 ;
		RECT 172.195 0.000 172.695 0.430 ;
		LAYER M2 ;
		RECT 194.290 0.000 194.790 0.430 ;
		LAYER VIA3 ;
		RECT 161.980 0.000 165.040 0.430 ;
		LAYER M3 ;
		RECT 161.980 0.000 165.040 0.430 ;
		LAYER M3 ;
		RECT 165.740 0.000 167.120 0.430 ;
		LAYER VIA3 ;
		RECT 165.740 0.000 167.120 0.430 ;
		LAYER M2 ;
		RECT 44.890 0.000 45.390 0.430 ;
		LAYER M3 ;
		RECT 34.690 0.000 35.790 0.430 ;
		LAYER M1 ;
		RECT 36.480 0.000 37.000 0.430 ;
		LAYER VIA3 ;
		RECT 44.890 0.000 45.390 0.430 ;
		LAYER VIA3 ;
		RECT 2.890 0.000 3.390 0.430 ;
		LAYER M1 ;
		RECT 2.880 0.000 3.400 0.430 ;
		LAYER M1 ;
		RECT 28.080 0.000 28.600 0.430 ;
		LAYER M2 ;
		RECT 28.090 0.000 28.590 0.430 ;
		LAYER M1 ;
		RECT 29.280 0.000 29.800 0.430 ;
		LAYER VIA3 ;
		RECT 34.690 0.000 35.790 0.430 ;
		LAYER VIA3 ;
		RECT 208.090 0.000 209.190 0.430 ;
		LAYER M1 ;
		RECT 203.880 0.000 205.000 0.430 ;
		LAYER M1 ;
		RECT 206.880 0.000 207.400 0.430 ;
		LAYER M2 ;
		RECT 206.890 0.000 207.390 0.430 ;
		LAYER M3 ;
		RECT 206.890 0.000 207.390 0.430 ;
		LAYER VIA3 ;
		RECT 206.890 0.000 207.390 0.430 ;
		LAYER M3 ;
		RECT 205.690 0.000 206.190 0.430 ;
		LAYER VIA3 ;
		RECT 205.690 0.000 206.190 0.430 ;
		LAYER M2 ;
		RECT 205.690 0.000 206.190 0.430 ;
		LAYER M1 ;
		RECT 205.680 0.000 206.200 0.430 ;
		LAYER M2 ;
		RECT 208.090 0.000 209.190 0.430 ;
		LAYER M2 ;
		RECT 202.690 0.000 203.190 0.430 ;
		LAYER M1 ;
		RECT 202.680 0.000 203.200 0.430 ;
		LAYER M1 ;
		RECT 199.680 0.000 200.800 0.430 ;
		LAYER M1 ;
		RECT 71.280 0.000 71.800 0.430 ;
		LAYER M3 ;
		RECT 71.290 0.000 71.790 0.430 ;
		LAYER VIA3 ;
		RECT 71.290 0.000 71.790 0.430 ;
		LAYER M2 ;
		RECT 71.290 0.000 71.790 0.430 ;
		LAYER VIA3 ;
		RECT 72.490 0.000 73.590 0.430 ;
		LAYER M2 ;
		RECT 72.490 0.000 73.590 0.430 ;
		LAYER M3 ;
		RECT 72.490 0.000 73.590 0.430 ;
		LAYER M3 ;
		RECT 74.290 0.000 74.790 0.430 ;
		LAYER M3 ;
		RECT 80.890 0.000 81.990 0.430 ;
		LAYER VIA3 ;
		RECT 80.890 0.000 81.990 0.430 ;
		LAYER M1 ;
		RECT 80.880 0.000 82.000 0.430 ;
		LAYER M1 ;
		RECT 83.880 0.000 84.400 0.430 ;
		LAYER M1 ;
		RECT 85.080 0.000 86.200 0.430 ;
		LAYER M3 ;
		RECT 86.890 0.000 87.390 0.430 ;
		LAYER M2 ;
		RECT 86.890 0.000 87.390 0.430 ;
		LAYER VIA3 ;
		RECT 74.290 0.000 74.790 0.430 ;
		LAYER M2 ;
		RECT 82.690 0.000 83.190 0.430 ;
		LAYER M3 ;
		RECT 82.690 0.000 83.190 0.430 ;
		LAYER M1 ;
		RECT 209.880 0.000 210.400 0.430 ;
		LAYER M2 ;
		RECT 215.290 0.000 215.790 0.430 ;
		LAYER M3 ;
		RECT 215.290 0.000 215.790 0.430 ;
		LAYER M1 ;
		RECT 211.080 0.000 211.600 0.430 ;
		LAYER VIA3 ;
		RECT 212.290 0.000 213.390 0.430 ;
		LAYER M2 ;
		RECT 214.090 0.000 214.590 0.430 ;
		LAYER M3 ;
		RECT 214.090 0.000 214.590 0.430 ;
		LAYER M1 ;
		RECT 158.210 0.000 161.290 0.430 ;
		LAYER M3 ;
		RECT 170.130 0.000 170.895 0.430 ;
		LAYER M1 ;
		RECT 165.730 0.000 167.130 0.430 ;
		LAYER M3 ;
		RECT 62.890 0.000 63.390 0.430 ;
		LAYER M3 ;
		RECT 61.690 0.000 62.190 0.430 ;
		LAYER M1 ;
		RECT 61.680 0.000 62.200 0.430 ;
		LAYER VIA3 ;
		RECT 64.090 0.000 65.190 0.430 ;
		LAYER M2 ;
		RECT 64.090 0.000 65.190 0.430 ;
		LAYER M2 ;
		RECT 65.890 0.000 66.390 0.430 ;
		LAYER M3 ;
		RECT 65.890 0.000 66.390 0.430 ;
		LAYER VIA3 ;
		RECT 65.890 0.000 66.390 0.430 ;
		LAYER M1 ;
		RECT 65.880 0.000 66.400 0.430 ;
		LAYER M2 ;
		RECT 67.090 0.000 67.590 0.430 ;
		LAYER M1 ;
		RECT 67.080 0.000 67.600 0.430 ;
		LAYER M1 ;
		RECT 64.080 0.000 65.200 0.430 ;
		LAYER VIA3 ;
		RECT 62.890 0.000 63.390 0.430 ;
		LAYER M2 ;
		RECT 62.890 0.000 63.390 0.430 ;
		LAYER VIA3 ;
		RECT 68.290 0.000 69.390 0.430 ;
		LAYER M3 ;
		RECT 44.890 0.000 45.390 0.430 ;
		LAYER M1 ;
		RECT 43.080 0.000 44.200 0.430 ;
		LAYER M2 ;
		RECT 40.690 0.000 41.190 0.430 ;
		LAYER M3 ;
		RECT 40.690 0.000 41.190 0.430 ;
		LAYER VIA3 ;
		RECT 40.690 0.000 41.190 0.430 ;
		LAYER M2 ;
		RECT 41.890 0.000 42.390 0.430 ;
		LAYER M2 ;
		RECT 2.890 0.000 3.390 0.430 ;
		LAYER M1 ;
		RECT 12.480 0.000 13.000 0.430 ;
		LAYER M1 ;
		RECT 8.280 0.000 8.800 0.430 ;
		LAYER VIA3 ;
		RECT 4.090 0.000 4.590 0.430 ;
		LAYER M1 ;
		RECT 5.280 0.000 6.400 0.430 ;
		LAYER M3 ;
		RECT 5.290 0.000 6.390 0.430 ;
		LAYER VIA3 ;
		RECT 5.290 0.000 6.390 0.430 ;
		LAYER VIA3 ;
		RECT 8.290 0.000 8.790 0.430 ;
		LAYER M2 ;
		RECT 5.290 0.000 6.390 0.430 ;
		LAYER M1 ;
		RECT 7.080 0.000 7.600 0.430 ;
		LAYER M3 ;
		RECT 7.090 0.000 7.590 0.430 ;
		LAYER VIA3 ;
		RECT 7.090 0.000 7.590 0.430 ;
		LAYER M3 ;
		RECT 8.290 0.000 8.790 0.430 ;
		LAYER M2 ;
		RECT 11.290 0.000 11.790 0.430 ;
		LAYER M1 ;
		RECT 9.480 0.000 10.600 0.430 ;
		LAYER M2 ;
		RECT 8.290 0.000 8.790 0.430 ;
		LAYER M2 ;
		RECT 13.690 0.000 14.790 0.430 ;
		LAYER M3 ;
		RECT 12.490 0.000 12.990 0.430 ;
		LAYER M3 ;
		RECT 46.090 0.000 46.590 0.430 ;
		LAYER M3 ;
		RECT 54.490 0.000 54.990 0.430 ;
		LAYER M3 ;
		RECT 55.690 0.000 56.790 0.430 ;
		LAYER VIA3 ;
		RECT 55.690 0.000 56.790 0.430 ;
		LAYER M1 ;
		RECT 44.880 0.000 45.400 0.430 ;
		LAYER VIA3 ;
		RECT 43.090 0.000 44.190 0.430 ;
		LAYER M3 ;
		RECT 41.890 0.000 42.390 0.430 ;
		LAYER M1 ;
		RECT 41.880 0.000 42.400 0.430 ;
		LAYER VIA3 ;
		RECT 46.090 0.000 46.590 0.430 ;
		LAYER M2 ;
		RECT 46.090 0.000 46.590 0.430 ;
		LAYER M3 ;
		RECT 2.890 0.000 3.390 0.430 ;
		LAYER M1 ;
		RECT 46.080 0.000 46.600 0.430 ;
		LAYER M2 ;
		RECT 53.290 0.000 53.790 0.430 ;
		LAYER M2 ;
		RECT 47.290 0.000 48.390 0.430 ;
		LAYER VIA3 ;
		RECT 47.290 0.000 48.390 0.430 ;
		LAYER M1 ;
		RECT 50.280 0.000 50.800 0.430 ;
		LAYER M2 ;
		RECT 51.490 0.000 52.590 0.430 ;
		LAYER M1 ;
		RECT 51.480 0.000 52.600 0.430 ;
		LAYER VIA3 ;
		RECT 53.290 0.000 53.790 0.430 ;
		LAYER M3 ;
		RECT 51.490 0.000 52.590 0.430 ;
		LAYER M3 ;
		RECT 53.290 0.000 53.790 0.430 ;
		LAYER M3 ;
		RECT 70.090 0.000 70.590 0.430 ;
		LAYER M2 ;
		RECT 70.090 0.000 70.590 0.430 ;
		LAYER M1 ;
		RECT 78.480 0.000 79.000 0.430 ;
		LAYER M1 ;
		RECT 72.480 0.000 73.600 0.430 ;
		LAYER M1 ;
		RECT 74.280 0.000 74.800 0.430 ;
		LAYER M2 ;
		RECT 78.490 0.000 78.990 0.430 ;
		LAYER M2 ;
		RECT 76.690 0.000 77.790 0.430 ;
		LAYER M3 ;
		RECT 76.690 0.000 77.790 0.430 ;
		LAYER VIA3 ;
		RECT 76.690 0.000 77.790 0.430 ;
		LAYER M3 ;
		RECT 75.490 0.000 75.990 0.430 ;
		LAYER M2 ;
		RECT 75.490 0.000 75.990 0.430 ;
		LAYER VIA3 ;
		RECT 75.490 0.000 75.990 0.430 ;
		LAYER M1 ;
		RECT 75.480 0.000 76.000 0.430 ;
		LAYER M3 ;
		RECT 78.490 0.000 78.990 0.430 ;
		LAYER VIA3 ;
		RECT 78.490 0.000 78.990 0.430 ;
		LAYER M2 ;
		RECT 74.290 0.000 74.790 0.430 ;
		LAYER M1 ;
		RECT 76.680 0.000 77.800 0.430 ;
		LAYER VIA3 ;
		RECT 32.290 0.000 32.790 0.430 ;
		LAYER M1 ;
		RECT 37.680 0.000 38.200 0.430 ;
		LAYER M3 ;
		RECT 38.890 0.000 39.990 0.430 ;
		LAYER M1 ;
		RECT 40.680 0.000 41.200 0.430 ;
		LAYER VIA3 ;
		RECT 38.890 0.000 39.990 0.430 ;
		LAYER M2 ;
		RECT 30.490 0.000 31.590 0.430 ;
		LAYER M2 ;
		RECT 9.490 0.000 10.590 0.430 ;
		LAYER M3 ;
		RECT 9.490 0.000 10.590 0.430 ;
		LAYER VIA3 ;
		RECT 9.490 0.000 10.590 0.430 ;
		LAYER M1 ;
		RECT 11.280 0.000 11.800 0.430 ;
		LAYER M3 ;
		RECT 11.290 0.000 11.790 0.430 ;
		LAYER VIA3 ;
		RECT 11.290 0.000 11.790 0.430 ;
		LAYER VIA3 ;
		RECT 12.490 0.000 12.990 0.430 ;
		LAYER M2 ;
		RECT 12.490 0.000 12.990 0.430 ;
		LAYER M3 ;
		RECT 22.090 0.000 23.190 0.430 ;
		LAYER M1 ;
		RECT 22.080 0.000 23.200 0.430 ;
		LAYER M1 ;
		RECT 13.680 0.000 14.800 0.430 ;
		LAYER M1 ;
		RECT 26.280 0.000 27.400 0.430 ;
		LAYER VIA3 ;
		RECT 23.890 0.000 24.390 0.430 ;
		LAYER M1 ;
		RECT 23.880 0.000 24.400 0.430 ;
		LAYER M1 ;
		RECT 25.080 0.000 25.600 0.430 ;
		LAYER M3 ;
		RECT 26.290 0.000 27.390 0.430 ;
		LAYER M2 ;
		RECT 25.090 0.000 25.590 0.430 ;
		LAYER M3 ;
		RECT 25.090 0.000 25.590 0.430 ;
		LAYER M2 ;
		RECT 23.890 0.000 24.390 0.430 ;
		LAYER M3 ;
		RECT 23.890 0.000 24.390 0.430 ;
		LAYER VIA3 ;
		RECT 25.090 0.000 25.590 0.430 ;
		LAYER VIA3 ;
		RECT 28.090 0.000 28.590 0.430 ;
		LAYER M3 ;
		RECT 28.090 0.000 28.590 0.430 ;
		LAYER M3 ;
		RECT 29.290 0.000 29.790 0.430 ;
		LAYER VIA3 ;
		RECT 29.290 0.000 29.790 0.430 ;
		LAYER VIA3 ;
		RECT 20.890 0.000 21.390 0.430 ;
		LAYER VIA3 ;
		RECT 19.690 0.000 20.190 0.430 ;
		LAYER M1 ;
		RECT 19.680 0.000 20.200 0.430 ;
		LAYER VIA3 ;
		RECT 13.690 0.000 14.790 0.430 ;
		LAYER VIA3 ;
		RECT 15.490 0.000 15.990 0.430 ;
		LAYER M3 ;
		RECT 15.490 0.000 15.990 0.430 ;
		LAYER M1 ;
		RECT 106.080 0.000 107.200 0.430 ;
		LAYER M2 ;
		RECT 106.090 0.000 107.190 0.430 ;
		LAYER VIA3 ;
		RECT 106.090 0.000 107.190 0.430 ;
		LAYER M2 ;
		RECT 113.290 0.000 113.790 0.430 ;
		LAYER VIA3 ;
		RECT 114.490 0.000 115.590 0.430 ;
		LAYER M1 ;
		RECT 114.480 0.000 115.600 0.430 ;
		LAYER M2 ;
		RECT 114.490 0.000 115.590 0.430 ;
		LAYER M3 ;
		RECT 114.490 0.000 115.590 0.430 ;
		LAYER VIA3 ;
		RECT 113.290 0.000 113.790 0.430 ;
		LAYER M2 ;
		RECT 116.290 0.000 116.790 0.430 ;
		LAYER M3 ;
		RECT 116.290 0.000 116.790 0.430 ;
		LAYER VIA3 ;
		RECT 116.290 0.000 116.790 0.430 ;
		LAYER M3 ;
		RECT 106.090 0.000 107.190 0.430 ;
		LAYER M2 ;
		RECT 110.290 0.000 111.390 0.430 ;
		LAYER M1 ;
		RECT 110.280 0.000 111.400 0.430 ;
		LAYER M3 ;
		RECT 110.290 0.000 111.390 0.430 ;
		LAYER VIA3 ;
		RECT 110.290 0.000 111.390 0.430 ;
		LAYER M3 ;
		RECT 107.890 0.000 108.390 0.430 ;
		LAYER M2 ;
		RECT 107.890 0.000 108.390 0.430 ;
		LAYER M1 ;
		RECT 109.080 0.000 109.600 0.430 ;
		LAYER M1 ;
		RECT 107.880 0.000 108.400 0.430 ;
		LAYER M2 ;
		RECT 109.090 0.000 109.590 0.430 ;
		LAYER M3 ;
		RECT 109.090 0.000 109.590 0.430 ;
		LAYER VIA3 ;
		RECT 109.090 0.000 109.590 0.430 ;
		LAYER VIA3 ;
		RECT 107.890 0.000 108.390 0.430 ;
		LAYER M1 ;
		RECT 113.280 0.000 113.800 0.430 ;
		LAYER M2 ;
		RECT 112.090 0.000 112.590 0.430 ;
		LAYER VIA3 ;
		RECT 112.090 0.000 112.590 0.430 ;
		LAYER M1 ;
		RECT 112.080 0.000 112.600 0.430 ;
		LAYER M3 ;
		RECT 113.290 0.000 113.790 0.430 ;
		LAYER M3 ;
		RECT 112.090 0.000 112.590 0.430 ;
		LAYER M2 ;
		RECT 97.690 0.000 98.790 0.430 ;
		LAYER VIA3 ;
		RECT 97.690 0.000 98.790 0.430 ;
		LAYER VIA3 ;
		RECT 99.490 0.000 99.990 0.430 ;
		LAYER VIA3 ;
		RECT 100.690 0.000 101.190 0.430 ;
		LAYER M2 ;
		RECT 158.220 0.000 161.280 0.430 ;
		LAYER VIA3 ;
		RECT 158.220 0.000 161.280 0.430 ;
		LAYER VIA3 ;
		RECT 103.690 0.000 104.190 0.430 ;
		LAYER M3 ;
		RECT 158.220 0.000 161.280 0.430 ;
		LAYER M1 ;
		RECT 103.680 0.000 104.200 0.430 ;
		LAYER M3 ;
		RECT 103.690 0.000 104.190 0.430 ;
		LAYER VIA3 ;
		RECT 101.890 0.000 102.990 0.430 ;
		LAYER M3 ;
		RECT 101.890 0.000 102.990 0.430 ;
		LAYER VIA3 ;
		RECT 104.890 0.000 105.390 0.430 ;
		LAYER M3 ;
		RECT 104.890 0.000 105.390 0.430 ;
		LAYER M1 ;
		RECT 104.880 0.000 105.400 0.430 ;
		LAYER M2 ;
		RECT 103.690 0.000 104.190 0.430 ;
		LAYER M2 ;
		RECT 104.890 0.000 105.390 0.430 ;
		LAYER M1 ;
		RECT 97.680 0.000 98.800 0.430 ;
		LAYER VIA3 ;
		RECT 95.290 0.000 95.790 0.430 ;
		LAYER M3 ;
		RECT 95.290 0.000 95.790 0.430 ;
		LAYER M3 ;
		RECT 100.690 0.000 101.190 0.430 ;
		LAYER M1 ;
		RECT 100.680 0.000 101.200 0.430 ;
		LAYER M2 ;
		RECT 99.490 0.000 99.990 0.430 ;
		LAYER M3 ;
		RECT 99.490 0.000 99.990 0.430 ;
		LAYER M2 ;
		RECT 100.690 0.000 101.190 0.430 ;
		LAYER M1 ;
		RECT 99.480 0.000 100.000 0.430 ;
		LAYER M1 ;
		RECT 101.880 0.000 103.000 0.430 ;
		LAYER M2 ;
		RECT 101.890 0.000 102.990 0.430 ;
		LAYER M3 ;
		RECT 97.690 0.000 98.790 0.430 ;
		LAYER M1 ;
		RECT 95.280 0.000 95.800 0.430 ;
		LAYER M2 ;
		RECT 95.290 0.000 95.790 0.430 ;
		LAYER M2 ;
		RECT 96.490 0.000 96.990 0.430 ;
		LAYER M3 ;
		RECT 96.490 0.000 96.990 0.430 ;
		LAYER VIA3 ;
		RECT 96.490 0.000 96.990 0.430 ;
		LAYER M1 ;
		RECT 96.480 0.000 97.000 0.430 ;
		LAYER M3 ;
		RECT 203.890 0.000 204.990 0.430 ;
		LAYER VIA3 ;
		RECT 202.690 0.000 203.190 0.430 ;
		LAYER M2 ;
		RECT 199.690 0.000 200.790 0.430 ;
		LAYER M1 ;
		RECT 201.480 0.000 202.000 0.430 ;
		LAYER M3 ;
		RECT 202.690 0.000 203.190 0.430 ;
		LAYER M2 ;
		RECT 201.490 0.000 201.990 0.430 ;
		LAYER M2 ;
		RECT 191.290 0.000 192.390 0.430 ;
		LAYER VIA3 ;
		RECT 191.290 0.000 192.390 0.430 ;
		LAYER M1 ;
		RECT 193.080 0.000 193.600 0.430 ;
		LAYER VIA3 ;
		RECT 201.490 0.000 201.990 0.430 ;
		LAYER M1 ;
		RECT 191.280 0.000 192.400 0.430 ;
		LAYER M3 ;
		RECT 191.290 0.000 192.390 0.430 ;
		LAYER M2 ;
		RECT 203.890 0.000 204.990 0.430 ;
		LAYER VIA3 ;
		RECT 203.890 0.000 204.990 0.430 ;
		LAYER VIA3 ;
		RECT 199.690 0.000 200.790 0.430 ;
		LAYER M3 ;
		RECT 176.445 0.000 176.945 0.430 ;
		LAYER M2 ;
		RECT 176.445 0.000 176.945 0.430 ;
		LAYER M2 ;
		RECT 167.820 0.000 169.430 0.430 ;
		LAYER VIA3 ;
		RECT 167.820 0.000 169.430 0.430 ;
		LAYER M3 ;
		RECT 167.820 0.000 169.430 0.430 ;
		LAYER M1 ;
		RECT 167.810 0.000 169.440 0.430 ;
		LAYER M2 ;
		RECT 161.980 0.000 165.040 0.430 ;
		LAYER M3 ;
		RECT 177.645 0.000 178.465 0.430 ;
		LAYER M1 ;
		RECT 161.970 0.000 165.050 0.430 ;
		LAYER M2 ;
		RECT 165.740 0.000 167.120 0.430 ;
		LAYER M1 ;
		RECT 184.535 0.000 185.085 0.430 ;
		LAYER M2 ;
		RECT 184.545 0.000 185.075 0.430 ;
		LAYER VIA3 ;
		RECT 184.545 0.000 185.075 0.430 ;
		LAYER M3 ;
		RECT 184.545 0.000 185.075 0.430 ;
		LAYER M3 ;
		RECT 185.775 0.000 186.900 0.430 ;
		LAYER VIA3 ;
		RECT 185.775 0.000 186.900 0.430 ;
		LAYER M2 ;
		RECT 185.775 0.000 186.900 0.430 ;
		LAYER M1 ;
		RECT 185.765 0.000 186.910 0.430 ;
		LAYER M3 ;
		RECT 187.600 0.000 188.190 0.430 ;
		LAYER VIA3 ;
		RECT 187.600 0.000 188.190 0.430 ;
		LAYER M1 ;
		RECT 187.590 0.000 188.200 0.430 ;
		LAYER M2 ;
		RECT 187.600 0.000 188.190 0.430 ;
		LAYER M3 ;
		RECT 188.890 0.000 189.390 0.430 ;
		LAYER M2 ;
		RECT 190.090 0.000 190.590 0.430 ;
		LAYER M1 ;
		RECT 190.080 0.000 190.600 0.430 ;
		LAYER M3 ;
		RECT 190.090 0.000 190.590 0.430 ;
		LAYER VIA3 ;
		RECT 190.090 0.000 190.590 0.430 ;
		LAYER M1 ;
		RECT 188.880 0.000 189.400 0.430 ;
		LAYER M2 ;
		RECT 181.975 0.000 182.645 0.430 ;
		LAYER VIA3 ;
		RECT 181.975 0.000 182.645 0.430 ;
		LAYER M1 ;
		RECT 181.965 0.000 182.655 0.430 ;
		LAYER M2 ;
		RECT 188.890 0.000 189.390 0.430 ;
		LAYER VIA3 ;
		RECT 188.890 0.000 189.390 0.430 ;
		LAYER M3 ;
		RECT 181.975 0.000 182.645 0.430 ;
		LAYER M2 ;
		RECT 180.455 0.000 181.275 0.430 ;
		LAYER M1 ;
		RECT 180.445 0.000 181.285 0.430 ;
		LAYER M1 ;
		RECT 179.155 0.000 179.165 0.430 ;
		LAYER M2 ;
		RECT 177.645 0.000 178.465 0.430 ;
		LAYER M1 ;
		RECT 176.435 0.000 176.955 0.430 ;
		LAYER VIA3 ;
		RECT 176.445 0.000 176.945 0.430 ;
		LAYER VIA3 ;
		RECT 170.130 0.000 170.895 0.430 ;
		LAYER M1 ;
		RECT 173.985 0.000 174.505 0.430 ;
		LAYER VIA3 ;
		RECT 172.195 0.000 172.695 0.430 ;
		LAYER M2 ;
		RECT 172.195 0.000 172.695 0.430 ;
		LAYER M1 ;
		RECT 172.185 0.000 172.705 0.430 ;
		LAYER M2 ;
		RECT 170.130 0.000 170.895 0.430 ;
		LAYER VIA3 ;
		RECT 180.455 0.000 181.275 0.430 ;
		LAYER M1 ;
		RECT 177.635 0.000 178.475 0.430 ;
		LAYER VIA3 ;
		RECT 177.645 0.000 178.465 0.430 ;
		LAYER M3 ;
		RECT 199.690 0.000 200.790 0.430 ;
		LAYER M1 ;
		RECT 197.280 0.000 197.800 0.430 ;
		LAYER M3 ;
		RECT 197.290 0.000 197.790 0.430 ;
		LAYER M3 ;
		RECT 201.490 0.000 201.990 0.430 ;
		LAYER M2 ;
		RECT 195.490 0.000 196.590 0.430 ;
		LAYER VIA3 ;
		RECT 195.490 0.000 196.590 0.430 ;
		LAYER M3 ;
		RECT 195.490 0.000 196.590 0.430 ;
		LAYER M1 ;
		RECT 195.480 0.000 196.600 0.430 ;
		LAYER VIA3 ;
		RECT 193.090 0.000 193.590 0.430 ;
		LAYER M2 ;
		RECT 193.090 0.000 193.590 0.430 ;
		LAYER M3 ;
		RECT 194.290 0.000 194.790 0.430 ;
		LAYER VIA3 ;
		RECT 194.290 0.000 194.790 0.430 ;
		LAYER M1 ;
		RECT 194.280 0.000 194.800 0.430 ;
		LAYER M3 ;
		RECT 193.090 0.000 193.590 0.430 ;
		LAYER M2 ;
		RECT 198.490 0.000 198.990 0.430 ;
		LAYER VIA3 ;
		RECT 198.490 0.000 198.990 0.430 ;
		LAYER M1 ;
		RECT 198.480 0.000 199.000 0.430 ;
		LAYER VIA3 ;
		RECT 197.290 0.000 197.790 0.430 ;
		LAYER M3 ;
		RECT 235.090 0.000 235.590 0.430 ;
		LAYER M2 ;
		RECT 247.690 0.000 248.190 0.430 ;
		LAYER M3 ;
		RECT 247.690 0.000 248.190 0.430 ;
		LAYER VIA3 ;
		RECT 247.690 0.000 248.190 0.430 ;
		LAYER M2 ;
		RECT 257.290 0.000 257.790 0.430 ;
		LAYER VIA3 ;
		RECT 257.290 0.000 257.790 0.430 ;
		LAYER M3 ;
		RECT 257.290 0.000 257.790 0.430 ;
		LAYER M1 ;
		RECT 257.280 0.000 257.800 0.430 ;
		LAYER M2 ;
		RECT 260.290 0.000 260.790 0.430 ;
		LAYER M1 ;
		RECT 260.280 0.000 260.800 0.430 ;
		LAYER M2 ;
		RECT 261.490 0.000 261.990 0.430 ;
		LAYER VIA3 ;
		RECT 261.490 0.000 261.990 0.430 ;
		LAYER M1 ;
		RECT 235.080 0.000 235.600 0.430 ;
		LAYER M2 ;
		RECT 240.490 0.000 240.990 0.430 ;
		LAYER M1 ;
		RECT 240.480 0.000 241.000 0.430 ;
		LAYER VIA3 ;
		RECT 241.690 0.000 242.790 0.430 ;
		LAYER M2 ;
		RECT 258.490 0.000 259.590 0.430 ;
		LAYER M3 ;
		RECT 258.490 0.000 259.590 0.430 ;
		LAYER VIA3 ;
		RECT 258.490 0.000 259.590 0.430 ;
		LAYER M1 ;
		RECT 258.480 0.000 259.600 0.430 ;
		LAYER M3 ;
		RECT 260.290 0.000 260.790 0.430 ;
		LAYER VIA3 ;
		RECT 260.290 0.000 260.790 0.430 ;
		LAYER M3 ;
		RECT 261.490 0.000 261.990 0.430 ;
		LAYER M2 ;
		RECT 256.090 0.000 256.590 0.430 ;
		LAYER M1 ;
		RECT 251.880 0.000 252.400 0.430 ;
		LAYER M3 ;
		RECT 250.090 0.000 251.190 0.430 ;
		LAYER M3 ;
		RECT 256.090 0.000 256.590 0.430 ;
		LAYER VIA3 ;
		RECT 256.090 0.000 256.590 0.430 ;
		LAYER M1 ;
		RECT 248.880 0.000 249.400 0.430 ;
		LAYER M1 ;
		RECT 256.080 0.000 256.600 0.430 ;
		LAYER M2 ;
		RECT 251.890 0.000 252.390 0.430 ;
		LAYER M3 ;
		RECT 251.890 0.000 252.390 0.430 ;
		LAYER VIA3 ;
		RECT 251.890 0.000 252.390 0.430 ;
		LAYER M1 ;
		RECT 253.080 0.000 253.600 0.430 ;
		LAYER M1 ;
		RECT 254.280 0.000 255.400 0.430 ;
		LAYER M3 ;
		RECT 254.290 0.000 255.390 0.430 ;
		LAYER M2 ;
		RECT 254.290 0.000 255.390 0.430 ;
		LAYER M2 ;
		RECT 253.090 0.000 253.590 0.430 ;
		LAYER M3 ;
		RECT 253.090 0.000 253.590 0.430 ;
		LAYER VIA3 ;
		RECT 253.090 0.000 253.590 0.430 ;
		LAYER VIA3 ;
		RECT 254.290 0.000 255.390 0.430 ;
		LAYER M3 ;
		RECT 248.890 0.000 249.390 0.430 ;
		LAYER M2 ;
		RECT 248.890 0.000 249.390 0.430 ;
		LAYER VIA3 ;
		RECT 248.890 0.000 249.390 0.430 ;
		LAYER M2 ;
		RECT 250.090 0.000 251.190 0.430 ;
		LAYER VIA3 ;
		RECT 235.090 0.000 235.590 0.430 ;
		LAYER M1 ;
		RECT 237.480 0.000 238.600 0.430 ;
		LAYER M3 ;
		RECT 237.490 0.000 238.590 0.430 ;
		LAYER M2 ;
		RECT 235.090 0.000 235.590 0.430 ;
		LAYER M2 ;
		RECT 236.290 0.000 236.790 0.430 ;
		LAYER M3 ;
		RECT 236.290 0.000 236.790 0.430 ;
		LAYER M1 ;
		RECT 236.280 0.000 236.800 0.430 ;
		LAYER M2 ;
		RECT 237.490 0.000 238.590 0.430 ;
		LAYER VIA3 ;
		RECT 236.290 0.000 236.790 0.430 ;
		LAYER VIA3 ;
		RECT 237.490 0.000 238.590 0.430 ;
		LAYER M3 ;
		RECT 244.690 0.000 245.190 0.430 ;
		LAYER VIA3 ;
		RECT 244.690 0.000 245.190 0.430 ;
		LAYER VIA3 ;
		RECT 245.890 0.000 246.990 0.430 ;
		LAYER M1 ;
		RECT 244.680 0.000 245.200 0.430 ;
		LAYER VIA3 ;
		RECT 243.490 0.000 243.990 0.430 ;
		LAYER M2 ;
		RECT 245.890 0.000 246.990 0.430 ;
		LAYER M3 ;
		RECT 245.890 0.000 246.990 0.430 ;
		LAYER M2 ;
		RECT 243.490 0.000 243.990 0.430 ;
		LAYER M3 ;
		RECT 227.890 0.000 228.390 0.430 ;
		LAYER M3 ;
		RECT 229.090 0.000 230.190 0.430 ;
		LAYER VIA3 ;
		RECT 229.090 0.000 230.190 0.430 ;
		LAYER M1 ;
		RECT 229.080 0.000 230.200 0.430 ;
		LAYER M2 ;
		RECT 229.090 0.000 230.190 0.430 ;
		LAYER M1 ;
		RECT 232.080 0.000 232.600 0.430 ;
		LAYER M2 ;
		RECT 230.890 0.000 231.390 0.430 ;
		LAYER M3 ;
		RECT 230.890 0.000 231.390 0.430 ;
		LAYER VIA3 ;
		RECT 230.890 0.000 231.390 0.430 ;
		LAYER M2 ;
		RECT 262.690 0.000 263.790 0.430 ;
		LAYER M3 ;
		RECT 262.690 0.000 263.790 0.430 ;
		LAYER M1 ;
		RECT 245.880 0.000 247.000 0.430 ;
		LAYER VIA3 ;
		RECT 262.690 0.000 263.790 0.430 ;
		LAYER M1 ;
		RECT 262.680 0.000 263.800 0.430 ;
		LAYER VIA3 ;
		RECT 227.890 0.000 228.390 0.430 ;
		LAYER M2 ;
		RECT 227.890 0.000 228.390 0.430 ;
		LAYER M1 ;
		RECT 230.880 0.000 231.400 0.430 ;
		LAYER M1 ;
		RECT 265.680 0.000 266.200 0.430 ;
		LAYER M3 ;
		RECT 271.090 0.000 272.190 0.430 ;
		LAYER M1 ;
		RECT 268.680 0.000 269.200 0.430 ;
		LAYER M3 ;
		RECT 269.890 0.000 270.390 0.430 ;
		LAYER M1 ;
		RECT 266.880 0.000 268.000 0.430 ;
		LAYER VIA3 ;
		RECT 271.090 0.000 272.190 0.430 ;
		LAYER M2 ;
		RECT 266.890 0.000 267.990 0.430 ;
		LAYER M3 ;
		RECT 266.890 0.000 267.990 0.430 ;
		LAYER VIA3 ;
		RECT 266.890 0.000 267.990 0.430 ;
		LAYER M2 ;
		RECT 268.690 0.000 269.190 0.430 ;
		LAYER M3 ;
		RECT 268.690 0.000 269.190 0.430 ;
		LAYER VIA3 ;
		RECT 268.690 0.000 269.190 0.430 ;
		LAYER M2 ;
		RECT 264.490 0.000 264.990 0.430 ;
		LAYER M3 ;
		RECT 264.490 0.000 264.990 0.430 ;
		LAYER M2 ;
		RECT 271.090 0.000 272.190 0.430 ;
		LAYER M1 ;
		RECT 261.480 0.000 262.000 0.430 ;
		LAYER VIA3 ;
		RECT 250.090 0.000 251.190 0.430 ;
		LAYER M1 ;
		RECT 250.080 0.000 251.200 0.430 ;
		LAYER M1 ;
		RECT 247.680 0.000 248.200 0.430 ;
		LAYER VIA3 ;
		RECT 233.290 0.000 234.390 0.430 ;
		LAYER M2 ;
		RECT 244.690 0.000 245.190 0.430 ;
		LAYER M3 ;
		RECT 241.690 0.000 242.790 0.430 ;
		LAYER M1 ;
		RECT 241.680 0.000 242.800 0.430 ;
		LAYER M1 ;
		RECT 239.280 0.000 239.800 0.430 ;
		LAYER M3 ;
		RECT 239.290 0.000 239.790 0.430 ;
		LAYER M2 ;
		RECT 239.290 0.000 239.790 0.430 ;
		LAYER VIA3 ;
		RECT 239.290 0.000 239.790 0.430 ;
		LAYER M3 ;
		RECT 240.490 0.000 240.990 0.430 ;
		LAYER VIA3 ;
		RECT 240.490 0.000 240.990 0.430 ;
		LAYER M2 ;
		RECT 241.690 0.000 242.790 0.430 ;
		LAYER M2 ;
		RECT 232.090 0.000 232.590 0.430 ;
		LAYER M3 ;
		RECT 232.090 0.000 232.590 0.430 ;
		LAYER VIA3 ;
		RECT 232.090 0.000 232.590 0.430 ;
		LAYER M1 ;
		RECT 233.280 0.000 234.400 0.430 ;
		LAYER M2 ;
		RECT 233.290 0.000 234.390 0.430 ;
		LAYER M3 ;
		RECT 233.290 0.000 234.390 0.430 ;
		LAYER M2 ;
		RECT 223.690 0.000 224.190 0.430 ;
		LAYER VIA3 ;
		RECT 223.690 0.000 224.190 0.430 ;
		LAYER M3 ;
		RECT 223.690 0.000 224.190 0.430 ;
		LAYER M3 ;
		RECT 224.890 0.000 225.990 0.430 ;
		LAYER M1 ;
		RECT 279.480 0.000 280.600 0.430 ;
		LAYER M1 ;
		RECT 278.280 0.000 278.800 0.430 ;
		LAYER M1 ;
		RECT 243.480 0.000 244.000 0.430 ;
		LAYER M3 ;
		RECT 279.490 0.000 280.590 0.430 ;
		LAYER VIA3 ;
		RECT 279.490 0.000 280.590 0.430 ;
		LAYER M2 ;
		RECT 274.090 0.000 274.590 0.430 ;
		LAYER M1 ;
		RECT 275.280 0.000 276.400 0.430 ;
		LAYER M2 ;
		RECT 277.090 0.000 277.590 0.430 ;
		LAYER M1 ;
		RECT 277.080 0.000 277.600 0.430 ;
		LAYER VIA3 ;
		RECT 274.090 0.000 274.590 0.430 ;
		LAYER M3 ;
		RECT 274.090 0.000 274.590 0.430 ;
		LAYER M2 ;
		RECT 278.290 0.000 278.790 0.430 ;
		LAYER M3 ;
		RECT 278.290 0.000 278.790 0.430 ;
		LAYER M2 ;
		RECT 222.490 0.000 222.990 0.430 ;
		LAYER M1 ;
		RECT 222.480 0.000 223.000 0.430 ;
		LAYER M1 ;
		RECT 226.680 0.000 227.200 0.430 ;
		LAYER M1 ;
		RECT 227.880 0.000 228.400 0.430 ;
		LAYER M1 ;
		RECT 220.680 0.000 221.800 0.430 ;
		LAYER M2 ;
		RECT 220.690 0.000 221.790 0.430 ;
		LAYER M1 ;
		RECT 223.680 0.000 224.200 0.430 ;
		LAYER VIA3 ;
		RECT 224.890 0.000 225.990 0.430 ;
		LAYER M2 ;
		RECT 224.890 0.000 225.990 0.430 ;
		LAYER M2 ;
		RECT 226.690 0.000 227.190 0.430 ;
		LAYER M3 ;
		RECT 226.690 0.000 227.190 0.430 ;
		LAYER VIA3 ;
		RECT 226.690 0.000 227.190 0.430 ;
		LAYER M1 ;
		RECT 224.880 0.000 226.000 0.430 ;
		LAYER M2 ;
		RECT 272.890 0.000 273.390 0.430 ;
		LAYER M1 ;
		RECT 272.880 0.000 273.400 0.430 ;
		LAYER M2 ;
		RECT 275.290 0.000 276.390 0.430 ;
		LAYER VIA3 ;
		RECT 275.290 0.000 276.390 0.430 ;
		LAYER VIA3 ;
		RECT 272.890 0.000 273.390 0.430 ;
		LAYER M3 ;
		RECT 272.890 0.000 273.390 0.430 ;
		LAYER VIA3 ;
		RECT 278.290 0.000 278.790 0.430 ;
		LAYER M3 ;
		RECT 275.290 0.000 276.390 0.430 ;
		LAYER M3 ;
		RECT 277.090 0.000 277.590 0.430 ;
		LAYER M3 ;
		RECT 222.490 0.000 222.990 0.430 ;
		LAYER VIA3 ;
		RECT 222.490 0.000 222.990 0.430 ;
		LAYER M3 ;
		RECT 243.490 0.000 243.990 0.430 ;
		LAYER M1 ;
		RECT 49.080 0.000 49.600 0.430 ;
		LAYER M3 ;
		RECT 49.090 0.000 49.590 0.430 ;
		LAYER VIA3 ;
		RECT 49.090 0.000 49.590 0.430 ;
		LAYER M3 ;
		RECT 47.290 0.000 48.390 0.430 ;
		LAYER M1 ;
		RECT 47.280 0.000 48.400 0.430 ;
		LAYER VIA3 ;
		RECT 86.890 0.000 87.390 0.430 ;
		LAYER M2 ;
		RECT 91.090 0.000 91.590 0.430 ;
		LAYER M3 ;
		RECT 91.090 0.000 91.590 0.430 ;
		LAYER M2 ;
		RECT 93.490 0.000 94.590 0.430 ;
		LAYER M1 ;
		RECT 89.280 0.000 90.400 0.430 ;
		LAYER VIA3 ;
		RECT 91.090 0.000 91.590 0.430 ;
		LAYER VIA3 ;
		RECT 50.290 0.000 50.790 0.430 ;
		LAYER M3 ;
		RECT 50.290 0.000 50.790 0.430 ;
		LAYER M2 ;
		RECT 50.290 0.000 50.790 0.430 ;
		LAYER VIA3 ;
		RECT 51.490 0.000 52.590 0.430 ;
		LAYER M1 ;
		RECT 53.280 0.000 53.800 0.430 ;
		LAYER M2 ;
		RECT 54.490 0.000 54.990 0.430 ;
		LAYER VIA3 ;
		RECT 54.490 0.000 54.990 0.430 ;
		LAYER M1 ;
		RECT 55.680 0.000 56.800 0.430 ;
		LAYER VIA3 ;
		RECT 57.490 0.000 57.990 0.430 ;
		LAYER M1 ;
		RECT 57.480 0.000 58.000 0.430 ;
		LAYER VIA3 ;
		RECT 59.890 0.000 60.990 0.430 ;
		LAYER M2 ;
		RECT 59.890 0.000 60.990 0.430 ;
		LAYER VIA3 ;
		RECT 61.690 0.000 62.190 0.430 ;
		LAYER M1 ;
		RECT 58.680 0.000 59.200 0.430 ;
		LAYER VIA3 ;
		RECT 85.090 0.000 86.190 0.430 ;
		LAYER M2 ;
		RECT 80.890 0.000 81.990 0.430 ;
		LAYER M2 ;
		RECT 79.690 0.000 80.190 0.430 ;
		LAYER M3 ;
		RECT 79.690 0.000 80.190 0.430 ;
		LAYER VIA3 ;
		RECT 79.690 0.000 80.190 0.430 ;
		LAYER M1 ;
		RECT 79.680 0.000 80.200 0.430 ;
		LAYER M1 ;
		RECT 62.880 0.000 63.400 0.430 ;
		LAYER M2 ;
		RECT 83.890 0.000 84.390 0.430 ;
		LAYER VIA3 ;
		RECT 83.890 0.000 84.390 0.430 ;
		LAYER M3 ;
		RECT 83.890 0.000 84.390 0.430 ;
		LAYER M2 ;
		RECT 85.090 0.000 86.190 0.430 ;
		LAYER VIA3 ;
		RECT 82.690 0.000 83.190 0.430 ;
		LAYER M1 ;
		RECT 82.680 0.000 83.200 0.430 ;
		LAYER M3 ;
		RECT 85.090 0.000 86.190 0.430 ;
		LAYER M3 ;
		RECT 88.090 0.000 88.590 0.430 ;
		LAYER VIA3 ;
		RECT 88.090 0.000 88.590 0.430 ;
		LAYER M2 ;
		RECT 88.090 0.000 88.590 0.430 ;
		LAYER M1 ;
		RECT 88.080 0.000 88.600 0.430 ;
		LAYER M1 ;
		RECT 86.880 0.000 87.400 0.430 ;
		LAYER M3 ;
		RECT 89.290 0.000 90.390 0.430 ;
		LAYER VIA3 ;
		RECT 89.290 0.000 90.390 0.430 ;
		LAYER M1 ;
		RECT 4.080 0.000 4.600 0.430 ;
		LAYER M2 ;
		RECT 4.090 0.000 4.590 0.430 ;
		LAYER M3 ;
		RECT 4.090 0.000 4.590 0.430 ;
		LAYER M2 ;
		RECT 7.090 0.000 7.590 0.430 ;
		LAYER M2 ;
		RECT 22.090 0.000 23.190 0.430 ;
		LAYER M3 ;
		RECT 20.890 0.000 21.390 0.430 ;
		LAYER M1 ;
		RECT 20.880 0.000 21.400 0.430 ;
		LAYER M3 ;
		RECT 19.690 0.000 20.190 0.430 ;
		LAYER VIA3 ;
		RECT 22.090 0.000 23.190 0.430 ;
		LAYER M1 ;
		RECT 17.880 0.000 19.000 0.430 ;
		LAYER VIA3 ;
		RECT 17.890 0.000 18.990 0.430 ;
		LAYER M3 ;
		RECT 13.690 0.000 14.790 0.430 ;
		LAYER M2 ;
		RECT 26.290 0.000 27.390 0.430 ;
		LAYER VIA3 ;
		RECT 26.290 0.000 27.390 0.430 ;
	END
	# End of OBS

END TS1N65LPHSA1024X64M4F

END LIBRARY
